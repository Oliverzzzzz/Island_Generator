<?xml version="1.0" encoding="ISO-8859-1"?>
<!DOCTYPE svg PUBLIC '-//W3C//DTD SVG 1.0//EN'
          'http://www.w3.org/TR/2001/REC-SVG-20010904/DTD/svg10.dtd'>
<svg xmlns:xlink="http://www.w3.org/1999/xlink" style="fill-opacity:1; color-rendering:auto; color-interpolation:auto; text-rendering:auto; stroke:black; stroke-linecap:square; stroke-miterlimit:10; shape-rendering:auto; stroke-opacity:1; fill:black; stroke-dasharray:none; font-weight:normal; stroke-width:1; font-family:'Dialog'; font-style:normal; stroke-linejoin:miter; font-size:12px; stroke-dashoffset:0; image-rendering:auto;" width="1920" height="1080" xmlns="http://www.w3.org/2000/svg"
><!--Generated by the Batik Graphics2D SVG Generator--><defs id="genericDefs"
  /><g
  ><g style="stroke-width:0.2;"
    ><path style="fill:none;" d="M808.7 0 L768.1 0 L770.4 33.42 L790.42 45.49 L808.99 29.99 L808.7 0 Z"
      /><path d="M808.7 0 L768.1 0 L770.4 33.42 L790.42 45.49 L808.99 29.99 L808.7 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1875.21 637.64 L1920 638.8 L1920 700.6 L1871.98 704 L1860.4301 694.84 L1875.21 637.64 Z"
      /><path d="M1875.21 637.64 L1920 638.8 L1920 700.6 L1871.98 704 L1860.4301 694.84 L1875.21 637.64 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1580.85 163.09 L1560.88 185.1 L1562.77 202.96 L1595.8199 218.17 L1627.9399 194.15 L1620.17 172.24 L1580.85 163.09 Z"
      /><path d="M1580.85 163.09 L1560.88 185.1 L1562.77 202.96 L1595.8199 218.17 L1627.9399 194.15 L1620.17 172.24 L1580.85 163.09 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1493.74 118.14 L1472.63 124.56 L1468.5601 170.61 L1484.6 186.25 L1495.34 187.86 L1523.46 165.28 L1523.54 140.17 L1493.74 118.14 Z"
      /><path d="M1493.74 118.14 L1472.63 124.56 L1468.5601 170.61 L1484.6 186.25 L1495.34 187.86 L1523.46 165.28 L1523.54 140.17 L1493.74 118.14 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M587.95 243.66 L609.28 265.25 L602.07 282.65 L570.81 285.57 L562.23 269.05 L587.95 243.66 Z"
      /><path d="M587.95 243.66 L609.28 265.25 L602.07 282.65 L570.81 285.57 L562.23 269.05 L587.95 243.66 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M145.36 468.54 L166.66 515.86 L156.76 525.29 L154.7 525.13 L126.08 499.72 L138.65 468.73 L145.36 468.54 Z"
      /><path d="M145.36 468.54 L166.66 515.86 L156.76 525.29 L154.7 525.13 L126.08 499.72 L138.65 468.73 L145.36 468.54 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M775.58 103.82 L766.15 92.92 L734.9 109.46 L733.39 121.2 L763.11 141.46 L772.63 139.14 L775.58 103.82 Z"
      /><path d="M775.58 103.82 L766.15 92.92 L734.9 109.46 L733.39 121.2 L763.11 141.46 L772.63 139.14 L775.58 103.82 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M240.95 841.26 L281.04 842.75 L283.98 847.14 L269.44 896.61 L223.55 881.63 L240.95 841.26 Z"
      /><path d="M240.95 841.26 L281.04 842.75 L283.98 847.14 L269.44 896.61 L223.55 881.63 L240.95 841.26 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M771.09 263.35 L806.92 279.76 L806.88 300.97 L784.24 319.04 L755.29 308.93 L747.88 278.67 L749.06 275.39 L771.09 263.35 Z"
      /><path d="M771.09 263.35 L806.92 279.76 L806.88 300.97 L784.24 319.04 L755.29 308.93 L747.88 278.67 L749.06 275.39 L771.09 263.35 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M726.63 704.85 L716.54 737.73 L670.4 745.89 L665.14 738.08 L664.09 707.68 L698.45 689.56 L726.63 704.85 Z"
      /><path d="M726.63 704.85 L716.54 737.73 L670.4 745.89 L665.14 738.08 L664.09 707.68 L698.45 689.56 L726.63 704.85 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M430.58 434.5 L418.39 439.75 L409.91 473.91 L440.49 488.16 L458.9 475.46 L462.49 460.86 L430.58 434.5 Z"
      /><path d="M430.58 434.5 L418.39 439.75 L409.91 473.91 L440.49 488.16 L458.9 475.46 L462.49 460.86 L430.58 434.5 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1176.76 241.35 L1138.6801 265.9 L1155.96 288.74 L1189.92 291.1 L1191.83 290.07 L1196.38 259.35 L1176.76 241.35 Z"
      /><path d="M1176.76 241.35 L1138.6801 265.9 L1155.96 288.74 L1189.92 291.1 L1191.83 290.07 L1196.38 259.35 L1176.76 241.35 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1746.54 602.05 L1801.49 611.6 L1809.28 636.85 L1804.1 649.95 L1779.63 665.45 L1748.97 660.26 L1729.78 626.92 L1746.54 602.05 Z"
      /><path d="M1746.54 602.05 L1801.49 611.6 L1809.28 636.85 L1804.1 649.95 L1779.63 665.45 L1748.97 660.26 L1729.78 626.92 L1746.54 602.05 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M440.55 713.32 L413.76 752.58 L382.83 728.75 L415.93 690.01 L440.55 713.32 Z"
      /><path d="M440.55 713.32 L413.76 752.58 L382.83 728.75 L415.93 690.01 L440.55 713.32 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1247.26 284.42 L1269.62 298.37 L1274.03 318.52 L1257.58 339.88 L1240.74 339.55 L1222.29 322.28 L1220.04 304.43 L1247.26 284.42 Z"
      /><path d="M1247.26 284.42 L1269.62 298.37 L1274.03 318.52 L1257.58 339.88 L1240.74 339.55 L1222.29 322.28 L1220.04 304.43 L1247.26 284.42 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1625.61 287.58 L1601.25 305.47 L1599.84 322.16 L1635.22 346.48 L1640.74 344.49 L1659.8101 307.07 L1659.65 306.49 L1625.61 287.58 Z"
      /><path d="M1625.61 287.58 L1601.25 305.47 L1599.84 322.16 L1635.22 346.48 L1640.74 344.49 L1659.8101 307.07 L1659.65 306.49 L1625.61 287.58 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M895.3 0 L844.9 0 L848.55 34.88 L892.55 25.16 L895.3 0 Z"
      /><path d="M895.3 0 L844.9 0 L848.55 34.88 L892.55 25.16 L895.3 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1044.1 592.7 L1063.46 621.71 L1043.42 652.95 L1003.36 623.23 L1004.55 613.8 L1044.1 592.7 Z"
      /><path d="M1044.1 592.7 L1063.46 621.71 L1043.42 652.95 L1003.36 623.23 L1004.55 613.8 L1044.1 592.7 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1501.39 467.72 L1509.12 471.17 L1521.04 501.48 L1501.65 522.45 L1463.17 496.76 L1473.84 476.71 L1501.39 467.72 Z"
      /><path d="M1501.39 467.72 L1509.12 471.17 L1521.04 501.48 L1501.65 522.45 L1463.17 496.76 L1473.84 476.71 L1501.39 467.72 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M53.35 86.93 L40.4 117 L0 115.4 L0 59.6 L30.34 58.6 L53.35 86.93 Z"
      /><path d="M53.35 86.93 L40.4 117 L0 115.4 L0 59.6 L30.34 58.6 L53.35 86.93 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1313.46 782.43 L1340.03 790.17 L1346.76 812.98 L1317.04 839.46 L1315.73 838.9 L1294.11 799.68 L1297.38 787.42 L1313.46 782.43 Z"
      /><path d="M1313.46 782.43 L1340.03 790.17 L1346.76 812.98 L1317.04 839.46 L1315.73 838.9 L1294.11 799.68 L1297.38 787.42 L1313.46 782.43 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1482.8 338.56 L1480.24 362.57 L1459.1899 380.18 L1443.3199 370.82 L1430.17 326.46 L1452.89 310.4 L1482.8 338.56 Z"
      /><path d="M1482.8 338.56 L1480.24 362.57 L1459.1899 380.18 L1443.3199 370.82 L1430.17 326.46 L1452.89 310.4 L1482.8 338.56 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M670.31 1013.63 L690.73 1036.8 L686.41 1048.59 L652.1 1054.14 L643.02 1035.6899 L670.31 1013.63 Z"
      /><path d="M670.31 1013.63 L690.73 1036.8 L686.41 1048.59 L652.1 1054.14 L643.02 1035.6899 L670.31 1013.63 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1088.38 325.73 L1111.92 347.33 L1091.98 373.07 L1064.61 366.4 L1059.17 332.18 L1088.38 325.73 Z"
      /><path d="M1088.38 325.73 L1111.92 347.33 L1091.98 373.07 L1064.61 366.4 L1059.17 332.18 L1088.38 325.73 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1147.47 640.99 L1102.33 619.32 L1099.2 621.85 L1093.29 670.76 L1126.7 678.55 L1143.8199 667.87 L1147.47 640.99 Z"
      /><path d="M1147.47 640.99 L1102.33 619.32 L1099.2 621.85 L1093.29 670.76 L1126.7 678.55 L1143.8199 667.87 L1147.47 640.99 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M272.99 157.66 L231.25 157.86 L228.02 160.6 L233.12 200.09 L245.73 207.9 L277.01 197.21 L272.99 157.66 Z"
      /><path d="M272.99 157.66 L231.25 157.86 L228.02 160.6 L233.12 200.09 L245.73 207.9 L277.01 197.21 L272.99 157.66 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M813.9 707.14 L783.58 687.58 L757.95 703.32 L775.8 745.34 L816.53 728.79 L813.9 707.14 Z"
      /><path d="M813.9 707.14 L783.58 687.58 L757.95 703.32 L775.8 745.34 L816.53 728.79 L813.9 707.14 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M343.81 691.25 L315.31 692.92 L307.49 703.68 L310.76 729.02 L351.05 747.2 L368.32 727.8 L359.3 702.33 L343.81 691.25 Z"
      /><path d="M343.81 691.25 L315.31 692.92 L307.49 703.68 L310.76 729.02 L351.05 747.2 L368.32 727.8 L359.3 702.33 L343.81 691.25 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M145.99 841.22 L180.3 855.2 L185.49 868.11 L157.58 900.48 L136.4 896.44 L122.35 863.2 L145.99 841.22 Z"
      /><path d="M145.99 841.22 L180.3 855.2 L185.49 868.11 L157.58 900.48 L136.4 896.44 L122.35 863.2 L145.99 841.22 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M80.89 211.7 L111.83 234.5 L92.84 267.22 L54.22 261.12 L51.94 252.8 L70.28 215.32 L80.89 211.7 Z"
      /><path d="M80.89 211.7 L111.83 234.5 L92.84 267.22 L54.22 261.12 L51.94 252.8 L70.28 215.32 L80.89 211.7 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1424.1 1028.36 L1447.71 1032.67 L1450.9 1080 L1393.7 1080 L1392.4399 1050.62 L1424.1 1028.36 Z"
      /><path d="M1424.1 1028.36 L1447.71 1032.67 L1450.9 1080 L1393.7 1080 L1392.4399 1050.62 L1424.1 1028.36 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1576.27 697.03 L1584.08 647.84 L1542.27 649.24 L1540.0699 684.66 L1571.35 700.37 L1576.27 697.03 Z"
      /><path d="M1576.27 697.03 L1584.08 647.84 L1542.27 649.24 L1540.0699 684.66 L1571.35 700.37 L1576.27 697.03 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M158.3 0 L101.4 0 L101.48 32.57 L146.04 44.13 L158.3 0 Z"
      /><path d="M158.3 0 L101.4 0 L101.48 32.57 L146.04 44.13 L158.3 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1380.6899 515.7 L1341.6801 508.91 L1338.6 510.38 L1331.91 531.87 L1342.1801 559.61 L1378.96 569.67 L1381.9301 568.38 L1380.6899 515.7 Z"
      /><path d="M1380.6899 515.7 L1341.6801 508.91 L1338.6 510.38 L1331.91 531.87 L1342.1801 559.61 L1378.96 569.67 L1381.9301 568.38 L1380.6899 515.7 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1783.5699 839.97 L1809.0699 876.86 L1795.61 898.36 L1756.09 895.2 L1752.73 843.92 L1783.5699 839.97 Z"
      /><path d="M1783.5699 839.97 L1809.0699 876.86 L1795.61 898.36 L1756.09 895.2 L1752.73 843.92 L1783.5699 839.97 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M43.3 622.13 L28.16 653.1 L0 654.4 L0 602.6 L43.3 622.13 Z"
      /><path d="M43.3 622.13 L28.16 653.1 L0 654.4 L0 602.6 L43.3 622.13 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1170.48 685.41 L1143.8199 667.87 L1126.7 678.55 L1127.3199 720.01 L1134.58 725.7 L1168.42 712.26 L1170.48 685.41 Z"
      /><path d="M1170.48 685.41 L1143.8199 667.87 L1126.7 678.55 L1127.3199 720.01 L1134.58 725.7 L1168.42 712.26 L1170.48 685.41 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1065.25 231.04 L1034.0699 196.01 L1003.76 199.86 L998.56 227.28 L1022.73 251.74 L1063.83 239.39 L1065.25 231.04 Z"
      /><path d="M1065.25 231.04 L1034.0699 196.01 L1003.76 199.86 L998.56 227.28 L1022.73 251.74 L1063.83 239.39 L1065.25 231.04 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1862.74 897.73 L1830.8 872.28 L1809.0699 876.86 L1795.61 898.36 L1806.26 928.94 L1825.4 934.44 L1861.58 905.02 L1862.74 897.73 Z"
      /><path d="M1862.74 897.73 L1830.8 872.28 L1809.0699 876.86 L1795.61 898.36 L1806.26 928.94 L1825.4 934.44 L1861.58 905.02 L1862.74 897.73 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M312.53 608.53 L342.26 634.64 L306.74 662.91 L284.04 650.54 L280.97 629.96 L312.53 608.53 Z"
      /><path d="M312.53 608.53 L342.26 634.64 L306.74 662.91 L284.04 650.54 L280.97 629.96 L312.53 608.53 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M253.38 725.63 L225.8 733.01 L216.28 745.45 L218.83 756.49 L254.85 786.24 L262.44 785.3 L284.39 757.45 L253.38 725.63 Z"
      /><path d="M253.38 725.63 L225.8 733.01 L216.28 745.45 L218.83 756.49 L254.85 786.24 L262.44 785.3 L284.39 757.45 L253.38 725.63 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1595.08 781.59 L1575.05 822.53 L1615.3101 837.22 L1628.54 831.63 L1621.48 788.64 L1595.08 781.59 Z"
      /><path d="M1595.08 781.59 L1575.05 822.53 L1615.3101 837.22 L1628.54 831.63 L1621.48 788.64 L1595.08 781.59 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M885.38 311.33 L862.79 302.24 L836.76 318.2 L837.35 351.49 L865.75 361.73 L891.65 326.99 L885.38 311.33 Z"
      /><path d="M885.38 311.33 L862.79 302.24 L836.76 318.2 L837.35 351.49 L865.75 361.73 L891.65 326.99 L885.38 311.33 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1610.7 0 L1554 0 L1550.71 37.38 L1598.03 52.39 L1610.7 0 Z"
      /><path d="M1610.7 0 L1554 0 L1550.71 37.38 L1598.03 52.39 L1610.7 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M565.74 546.27 L578.67 553.44 L583.21 565.78 L575.39 590.19 L563.53 596.4 L550.84 594.4 L528.65 568.24 L528.58 567.54 L565.74 546.27 Z"
      /><path d="M565.74 546.27 L578.67 553.44 L583.21 565.78 L575.39 590.19 L563.53 596.4 L550.84 594.4 L528.65 568.24 L528.58 567.54 L565.74 546.27 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M494.34 229.32 L450.27 232.61 L453.65 266.38 L480.97 274.71 L495.02 261.75 L494.34 229.32 Z"
      /><path d="M494.34 229.32 L450.27 232.61 L453.65 266.38 L480.97 274.71 L495.02 261.75 L494.34 229.32 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1084.63 923.49 L1067.77 922.53 L1041.51 949 L1057.75 975.91 L1070.26 977.26 L1092.38 944.08 L1084.63 923.49 Z"
      /><path d="M1084.63 923.49 L1067.77 922.53 L1041.51 949 L1057.75 975.91 L1070.26 977.26 L1092.38 944.08 L1084.63 923.49 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1635.22 346.48 L1599.84 322.16 L1578.22 340.14 L1576.6801 351.18 L1609.1801 379.36 L1617.1801 380.46 L1635.22 346.48 Z"
      /><path d="M1635.22 346.48 L1599.84 322.16 L1578.22 340.14 L1576.6801 351.18 L1609.1801 379.36 L1617.1801 380.46 L1635.22 346.48 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1482.29 56.07 L1455.37 59.71 L1455.34 59.75 L1448.14 100.48 L1457.83 117.45 L1472.63 124.56 L1493.74 118.14 L1505.4301 86.27 L1482.29 56.07 Z"
      /><path d="M1482.29 56.07 L1455.37 59.71 L1455.34 59.75 L1448.14 100.48 L1457.83 117.45 L1472.63 124.56 L1493.74 118.14 L1505.4301 86.27 L1482.29 56.07 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M634.66 239.16 L665.99 255.76 L650.41 287.31 L622.21 261.34 L634.66 239.16 Z"
      /><path d="M634.66 239.16 L665.99 255.76 L650.41 287.31 L622.21 261.34 L634.66 239.16 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1920 287.1 L1920 347.8 L1887.2 345.36 L1878.89 291.32 L1920 287.1 Z"
      /><path d="M1920 287.1 L1920 347.8 L1887.2 345.36 L1878.89 291.32 L1920 287.1 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1226.0699 115.48 L1192.15 145.76 L1192.65 164.59 L1199.71 173.23 L1247.72 167.9 L1254.64 141.09 L1249.65 129.63 L1226.0699 115.48 Z"
      /><path d="M1226.0699 115.48 L1192.15 145.76 L1192.65 164.59 L1199.71 173.23 L1247.72 167.9 L1254.64 141.09 L1249.65 129.63 L1226.0699 115.48 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M746.88 165.35 L750.89 180.08 L740.8 191.59 L715.04 191.51 L702.6 176.55 L721.54 155.66 L746.88 165.35 Z"
      /><path d="M746.88 165.35 L750.89 180.08 L740.8 191.59 L715.04 191.51 L702.6 176.55 L721.54 155.66 L746.88 165.35 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M733.03 329.54 L731.27 352.79 L679.89 348.47 L677.02 341.68 L700.69 307.47 L733.03 329.54 Z"
      /><path d="M733.03 329.54 L731.27 352.79 L679.89 348.47 L677.02 341.68 L700.69 307.47 L733.03 329.54 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M408.31 840.08 L415.5 841.26 L442.61 882.65 L440 896.48 L432.29 904.38 L400.96 910.48 L374.42 881.95 L377.79 862.57 L408.31 840.08 Z"
      /><path d="M408.31 840.08 L415.5 841.26 L442.61 882.65 L440 896.48 L432.29 904.38 L400.96 910.48 L374.42 881.95 L377.79 862.57 L408.31 840.08 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M615.81 984.44 L633.99 989.74 L628.58 1029.45 L605.81 1036.52 L601.86 1034.64 L590.03 996.39 L590.69 995.21 L615.81 984.44 Z"
      /><path d="M615.81 984.44 L633.99 989.74 L628.58 1029.45 L605.81 1036.52 L601.86 1034.64 L590.03 996.39 L590.69 995.21 L615.81 984.44 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M837.35 351.49 L865.75 361.73 L873.69 377.34 L859.8 411.53 L819.78 407.99 L817.05 364.42 L837.35 351.49 Z"
      /><path d="M837.35 351.49 L865.75 361.73 L873.69 377.34 L859.8 411.53 L819.78 407.99 L817.05 364.42 L837.35 351.49 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M578.64 45.89 L562.5 33.46 L527.47 47.56 L527.64 70.85 L550.41 85.84 L577.13 72.25 L578.64 45.89 Z"
      /><path d="M578.64 45.89 L562.5 33.46 L527.47 47.56 L527.64 70.85 L550.41 85.84 L577.13 72.25 L578.64 45.89 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M0 816.6 L44.8 827.22 L51.24 843.16 L34.29 872.34 L0 874 L0 816.6 Z"
      /><path d="M0 816.6 L44.8 827.22 L51.24 843.16 L34.29 872.34 L0 874 L0 816.6 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1853.9399 68.19 L1856.04 69.2 L1875.45 105.09 L1870.74 118.59 L1849.27 127.73 L1821.16 109.76 L1839.3101 70.88 L1853.9399 68.19 Z"
      /><path d="M1853.9399 68.19 L1856.04 69.2 L1875.45 105.09 L1870.74 118.59 L1849.27 127.73 L1821.16 109.76 L1839.3101 70.88 L1853.9399 68.19 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1538.33 79.6 L1555.86 96.13 L1559.1899 119.08 L1523.54 140.17 L1493.74 118.14 L1505.4301 86.27 L1538.33 79.6 Z"
      /><path d="M1538.33 79.6 L1555.86 96.13 L1559.1899 119.08 L1523.54 140.17 L1493.74 118.14 L1505.4301 86.27 L1538.33 79.6 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1517.8 387.69 L1494.58 416.59 L1494.96 423.23 L1533.52 431.66 L1544.29 403.91 L1517.8 387.69 Z"
      /><path d="M1517.8 387.69 L1494.58 416.59 L1494.96 423.23 L1533.52 431.66 L1544.29 403.91 L1517.8 387.69 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1920 473.8 L1920 494.1 L1858.72 507.52 L1842.1899 459.25 L1857.52 440.85 L1866.89 439.35 L1920 473.8 Z"
      /><path d="M1920 473.8 L1920 494.1 L1858.72 507.52 L1842.1899 459.25 L1857.52 440.85 L1866.89 439.35 L1920 473.8 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M522.86 790.57 L515.71 781.42 L460.19 811.18 L488.41 851.34 L513.68 839.55 L522.86 790.57 Z"
      /><path d="M522.86 790.57 L515.71 781.42 L460.19 811.18 L488.41 851.34 L513.68 839.55 L522.86 790.57 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1557.05 263.13 L1565.6899 268.2 L1569.16 282.21 L1546.6801 316.56 L1523.41 320.71 L1521.74 319.76 L1513.58 300.32 L1526.48 269.61 L1557.05 263.13 Z"
      /><path d="M1557.05 263.13 L1565.6899 268.2 L1569.16 282.21 L1546.6801 316.56 L1523.41 320.71 L1521.74 319.76 L1513.58 300.32 L1526.48 269.61 L1557.05 263.13 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M185.49 868.11 L220.47 883.01 L211.35 923.47 L175.39 935 L157.58 900.48 L185.49 868.11 Z"
      /><path d="M185.49 868.11 L220.47 883.01 L211.35 923.47 L175.39 935 L157.58 900.48 L185.49 868.11 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1472.63 124.56 L1457.83 117.45 L1418.35 145.5 L1426.51 174.53 L1468.5601 170.61 L1472.63 124.56 Z"
      /><path d="M1472.63 124.56 L1457.83 117.45 L1418.35 145.5 L1426.51 174.53 L1468.5601 170.61 L1472.63 124.56 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1742.8 376.59 L1703.4399 332.07 L1676.96 366.67 L1680.42 390 L1742.84 378.24 L1742.8 376.59 Z"
      /><path d="M1742.8 376.59 L1703.4399 332.07 L1676.96 366.67 L1680.42 390 L1742.84 378.24 L1742.8 376.59 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M852.39 1009.18 L820.08 1029.89 L818.2 1080 L869.8 1080 L866.53 1022.19 L856.7 1011.05 L852.39 1009.18 Z"
      /><path d="M852.39 1009.18 L820.08 1029.89 L818.2 1080 L869.8 1080 L866.53 1022.19 L856.7 1011.05 L852.39 1009.18 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1920 841.1 L1920 799 L1867.73 802.62 L1857.02 826.37 L1883.42 848.34 L1920 841.1 Z"
      /><path d="M1920 841.1 L1920 799 L1867.73 802.62 L1857.02 826.37 L1883.42 848.34 L1920 841.1 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1468.5601 170.61 L1484.6 186.25 L1450.51 231.38 L1439.97 232.47 L1433.16 226.39 L1426.0699 175.24 L1426.51 174.53 L1468.5601 170.61 Z"
      /><path d="M1468.5601 170.61 L1484.6 186.25 L1450.51 231.38 L1439.97 232.47 L1433.16 226.39 L1426.0699 175.24 L1426.51 174.53 L1468.5601 170.61 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1634.17 1041.53 L1665.23 1063.58 L1666.2 1080 L1609.1 1080 L1613.15 1052.92 L1634.17 1041.53 Z"
      /><path d="M1634.17 1041.53 L1665.23 1063.58 L1666.2 1080 L1609.1 1080 L1613.15 1052.92 L1634.17 1041.53 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M684.44 928.07 L649.86 919.29 L634.69 937.7 L650.15 961.81 L678.49 962.32 L688.12 950.21 L684.44 928.07 Z"
      /><path d="M684.44 928.07 L649.86 919.29 L634.69 937.7 L650.15 961.81 L678.49 962.32 L688.12 950.21 L684.44 928.07 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M526.08 273.91 L495.02 261.75 L480.97 274.71 L484.25 299.79 L522.95 305.37 L526.08 273.91 Z"
      /><path d="M526.08 273.91 L495.02 261.75 L480.97 274.71 L484.25 299.79 L522.95 305.37 L526.08 273.91 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M780.35 187.15 L813.92 198.14 L819.05 213.36 L807.56 229.46 L776.4 231.33 L771.31 225.5 L778.92 187.9 L780.35 187.15 Z"
      /><path d="M780.35 187.15 L813.92 198.14 L819.05 213.36 L807.56 229.46 L776.4 231.33 L771.31 225.5 L778.92 187.9 L780.35 187.15 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1192.65 164.59 L1143.4 177.01 L1143.95 206.5 L1175.3199 222.58 L1200.14 201.37 L1199.71 173.23 L1192.65 164.59 Z"
      /><path d="M1192.65 164.59 L1143.4 177.01 L1143.95 206.5 L1175.3199 222.58 L1200.14 201.37 L1199.71 173.23 L1192.65 164.59 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1813.6801 525.98 L1801.72 558.53 L1754.4301 557.35 L1760.46 508.52 L1791.53 503.05 L1813.6801 525.98 Z"
      /><path d="M1813.6801 525.98 L1801.72 558.53 L1754.4301 557.35 L1760.46 508.52 L1791.53 503.05 L1813.6801 525.98 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M838.49 573.12 L795.53 574.95 L791.61 578.53 L795.29 610.68 L824.03 628.74 L845.64 618.62 L852.86 597.26 L838.49 573.12 Z"
      /><path d="M838.49 573.12 L795.53 574.95 L791.61 578.53 L795.29 610.68 L824.03 628.74 L845.64 618.62 L852.86 597.26 L838.49 573.12 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M731.27 1031.6801 L728 1080 L698.2 1080 L686.41 1048.59 L690.73 1036.8 L720.88 1024.34 L731.27 1031.6801 Z"
      /><path d="M731.27 1031.6801 L728 1080 L698.2 1080 L686.41 1048.59 L690.73 1036.8 L720.88 1024.34 L731.27 1031.6801 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M778.44 511.21 L798.01 524.54 L795.53 574.95 L791.61 578.53 L764.33 575.07 L746.84 543.03 L769.17 513.28 L778.44 511.21 Z"
      /><path d="M778.44 511.21 L798.01 524.54 L795.53 574.95 L791.61 578.53 L764.33 575.07 L746.84 543.03 L769.17 513.28 L778.44 511.21 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M221.03 494.45 L205.17 530.29 L175.66 513.11 L187.54 491.78 L214.8 486.24 L221.03 494.45 Z"
      /><path d="M221.03 494.45 L205.17 530.29 L175.66 513.11 L187.54 491.78 L214.8 486.24 L221.03 494.45 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1438.49 421.87 L1444.3101 437.91 L1425.3101 457.51 L1382.34 447.77 L1396.95 405.91 L1438.49 421.87 Z"
      /><path d="M1438.49 421.87 L1444.3101 437.91 L1425.3101 457.51 L1382.34 447.77 L1396.95 405.91 L1438.49 421.87 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1342.1 736.29 L1356 772.05 L1340.03 790.17 L1313.46 782.43 L1326.7 732.88 L1327.24 732.39 L1342.1 736.29 Z"
      /><path d="M1342.1 736.29 L1356 772.05 L1340.03 790.17 L1313.46 782.43 L1326.7 732.88 L1327.24 732.39 L1342.1 736.29 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M686.41 1048.59 L652.1 1054.14 L644.6 1080 L698.2 1080 L686.41 1048.59 Z"
      /><path d="M686.41 1048.59 L652.1 1054.14 L644.6 1080 L698.2 1080 L686.41 1048.59 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M550.84 594.4 L528.65 568.24 L498.36 605.97 L501.58 621.08 L529.66 623 L550.84 594.4 Z"
      /><path d="M550.84 594.4 L528.65 568.24 L498.36 605.97 L501.58 621.08 L529.66 623 L550.84 594.4 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M340.74 376.24 L308.51 369.58 L288.51 396.82 L331.64 418.05 L346.18 392.15 L340.74 376.24 Z"
      /><path d="M340.74 376.24 L308.51 369.58 L288.51 396.82 L331.64 418.05 L346.18 392.15 L340.74 376.24 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1721.23 700.74 L1677.38 663.45 L1671.25 664.74 L1656.27 706.76 L1696.33 732.66 L1721.49 704.34 L1721.23 700.74 Z"
      /><path d="M1721.23 700.74 L1677.38 663.45 L1671.25 664.74 L1656.27 706.76 L1696.33 732.66 L1721.49 704.34 L1721.23 700.74 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M450.27 232.61 L442.9 226.34 L402.77 250.57 L414.86 281.7 L425.82 285.88 L433.6 284.63 L453.65 266.38 L450.27 232.61 Z"
      /><path d="M450.27 232.61 L442.9 226.34 L402.77 250.57 L414.86 281.7 L425.82 285.88 L433.6 284.63 L453.65 266.38 L450.27 232.61 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M908.74 529.58 L939.23 541.11 L947.93 587.73 L938.81 598.18 L905.57 599.27 L894.65 590.01 L893.09 546.65 L908.74 529.58 Z"
      /><path d="M908.74 529.58 L939.23 541.11 L947.93 587.73 L938.81 598.18 L905.57 599.27 L894.65 590.01 L893.09 546.65 L908.74 529.58 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M38.41 559.12 L0.92 537.07 L0 537.1 L0 593.4 L37.53 573.98 L38.41 559.12 Z"
      /><path d="M38.41 559.12 L0.92 537.07 L0 537.1 L0 593.4 L37.53 573.98 L38.41 559.12 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1379.4399 685.11 L1418.3101 716.35 L1417.35 737.13 L1398.35 750.09 L1366.34 725.41 L1379.4399 685.11 Z"
      /><path d="M1379.4399 685.11 L1418.3101 716.35 L1417.35 737.13 L1398.35 750.09 L1366.34 725.41 L1379.4399 685.11 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M626.47 76.3 L644.65 89.57 L647.01 119.64 L595.02 127.31 L594.41 126.09 L599.39 87.83 L626.47 76.3 Z"
      /><path d="M626.47 76.3 L644.65 89.57 L647.01 119.64 L595.02 127.31 L594.41 126.09 L599.39 87.83 L626.47 76.3 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M683.86 608.36 L669.14 610 L661.32 616.96 L658.71 648.64 L661.1 653.16 L694.49 657.67 L704.99 646.62 L701.91 621.12 L683.86 608.36 Z"
      /><path d="M683.86 608.36 L669.14 610 L661.32 616.96 L658.71 648.64 L661.1 653.16 L694.49 657.67 L704.99 646.62 L701.91 621.12 L683.86 608.36 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M740.09 652.32 L704.99 646.62 L694.49 657.67 L698.45 689.56 L726.63 704.85 L739.87 699.1 L740.09 652.32 Z"
      /><path d="M740.09 652.32 L704.99 646.62 L694.49 657.67 L698.45 689.56 L726.63 704.85 L739.87 699.1 L740.09 652.32 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M959.39 135.15 L957 136.4 L955.41 186.63 L999.01 194.34 L1001.79 146.38 L959.39 135.15 Z"
      /><path d="M959.39 135.15 L957 136.4 L955.41 186.63 L999.01 194.34 L1001.79 146.38 L959.39 135.15 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M355.54 287.5 L346.14 290.12 L320.97 323.75 L320.99 324.12 L354.79 348.54 L358.13 347.46 L374.39 301.88 L355.54 287.5 Z"
      /><path d="M355.54 287.5 L346.14 290.12 L320.97 323.75 L320.99 324.12 L354.79 348.54 L358.13 347.46 L374.39 301.88 L355.54 287.5 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1570.7 923.06 L1580.21 964.78 L1563.1801 975.38 L1519.88 964.62 L1524.03 932.1 L1559.99 917.44 L1570.7 923.06 Z"
      /><path d="M1570.7 923.06 L1580.21 964.78 L1563.1801 975.38 L1519.88 964.62 L1524.03 932.1 L1559.99 917.44 L1570.7 923.06 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M884.22 69.05 L897.16 101.89 L869.37 120.26 L847.11 96.01 L855.28 66.81 L884.22 69.05 Z"
      /><path d="M884.22 69.05 L897.16 101.89 L869.37 120.26 L847.11 96.01 L855.28 66.81 L884.22 69.05 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M159.68 762.89 L156.91 761.78 L125.76 773.69 L119.69 804.35 L141.94 817.71 L173.24 794.54 L159.68 762.89 Z"
      /><path d="M159.68 762.89 L156.91 761.78 L125.76 773.69 L119.69 804.35 L141.94 817.71 L173.24 794.54 L159.68 762.89 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1604.86 65.37 L1614.66 71.38 L1607.83 117.67 L1575.74 129.81 L1559.1899 119.08 L1555.86 96.13 L1604.86 65.37 Z"
      /><path d="M1604.86 65.37 L1614.66 71.38 L1607.83 117.67 L1575.74 129.81 L1559.1899 119.08 L1555.86 96.13 L1604.86 65.37 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M354.28 521.07 L379.05 526.24 L386.89 567.06 L359.64 580.4 L342.17 573.17 L332.53 537.24 L354.28 521.07 Z"
      /><path d="M354.28 521.07 L379.05 526.24 L386.89 567.06 L359.64 580.4 L342.17 573.17 L332.53 537.24 L354.28 521.07 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1443.3199 370.82 L1398.83 382.64 L1392.42 393.75 L1396.95 405.91 L1438.49 421.87 L1459.28 381.03 L1459.1899 380.18 L1443.3199 370.82 Z"
      /><path d="M1443.3199 370.82 L1398.83 382.64 L1392.42 393.75 L1396.95 405.91 L1438.49 421.87 L1459.28 381.03 L1459.1899 380.18 L1443.3199 370.82 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M196.63 340.12 L184.49 333.54 L143.75 349.94 L158.05 393.14 L192.2 387.02 L196.63 340.12 Z"
      /><path d="M196.63 340.12 L184.49 333.54 L143.75 349.94 L158.05 393.14 L192.2 387.02 L196.63 340.12 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1607.67 519.21 L1585.85 512.55 L1562.9399 523.64 L1560.25 538.15 L1592.5 568.56 L1610.71 565.86 L1622.1801 548.17 L1607.67 519.21 Z"
      /><path d="M1607.67 519.21 L1585.85 512.55 L1562.9399 523.64 L1560.25 538.15 L1592.5 568.56 L1610.71 565.86 L1622.1801 548.17 L1607.67 519.21 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1499.6899 907.95 L1478.34 909.48 L1462.87 928.99 L1486.05 973.14 L1509.52 973.32 L1519.88 964.62 L1524.03 932.1 L1499.6899 907.95 Z"
      /><path d="M1499.6899 907.95 L1478.34 909.48 L1462.87 928.99 L1486.05 973.14 L1509.52 973.32 L1519.88 964.62 L1524.03 932.1 L1499.6899 907.95 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M216.25 569.85 L241.26 569.85 L249.23 583.1 L216.99 614.51 L204.59 599.81 L216.25 569.85 Z"
      /><path d="M216.25 569.85 L241.26 569.85 L249.23 583.1 L216.99 614.51 L204.59 599.81 L216.25 569.85 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1059.17 332.18 L1058.8101 331.92 L1022.96 332.49 L1021.63 383.02 L1040.53 386.28 L1064.61 366.4 L1059.17 332.18 Z"
      /><path d="M1059.17 332.18 L1058.8101 331.92 L1022.96 332.49 L1021.63 383.02 L1040.53 386.28 L1064.61 366.4 L1059.17 332.18 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1376.49 451.74 L1396.39 505.84 L1380.6899 515.7 L1341.6801 508.91 L1356.74 452.47 L1376.49 451.74 Z"
      /><path d="M1376.49 451.74 L1396.39 505.84 L1380.6899 515.7 L1341.6801 508.91 L1356.74 452.47 L1376.49 451.74 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M323.82 89.61 L347.01 113.6 L329.63 145.78 L328.7 145.89 L301.14 106.97 L301.85 103.1 L323.82 89.61 Z"
      /><path d="M323.82 89.61 L347.01 113.6 L329.63 145.78 L328.7 145.89 L301.14 106.97 L301.85 103.1 L323.82 89.61 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1428.72 265.91 L1385.4301 280.58 L1419.4399 325.79 L1430.17 326.46 L1452.89 310.4 L1455.78 299.92 L1428.72 265.91 Z"
      /><path d="M1428.72 265.91 L1385.4301 280.58 L1419.4399 325.79 L1430.17 326.46 L1452.89 310.4 L1455.78 299.92 L1428.72 265.91 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M845.28 54.12 L855.28 66.81 L847.11 96.01 L816.09 102.58 L809.08 71.91 L845.28 54.12 Z"
      /><path d="M845.28 54.12 L855.28 66.81 L847.11 96.01 L816.09 102.58 L809.08 71.91 L845.28 54.12 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M386.27 398.57 L388.43 423.74 L364.5 444.16 L332.83 426.99 L331.64 418.05 L346.18 392.15 L386.27 398.57 Z"
      /><path d="M386.27 398.57 L388.43 423.74 L364.5 444.16 L332.83 426.99 L331.64 418.05 L346.18 392.15 L386.27 398.57 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1185.5699 413.55 L1160.48 442.07 L1171.85 469.55 L1209.3199 465.89 L1220.26 440.25 L1201.66 415.02 L1185.5699 413.55 Z"
      /><path d="M1185.5699 413.55 L1160.48 442.07 L1171.85 469.55 L1209.3199 465.89 L1220.26 440.25 L1201.66 415.02 L1185.5699 413.55 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M374.04 110.31 L347.01 113.6 L323.82 89.61 L328.15 78.14 L371 73.63 L374.04 110.31 Z"
      /><path d="M374.04 110.31 L347.01 113.6 L323.82 89.61 L328.15 78.14 L371 73.63 L374.04 110.31 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1259.36 186.73 L1257.5699 201.83 L1230.11 220.28 L1200.14 201.37 L1199.71 173.23 L1247.72 167.9 L1259.36 186.73 Z"
      /><path d="M1259.36 186.73 L1257.5699 201.83 L1230.11 220.28 L1200.14 201.37 L1199.71 173.23 L1247.72 167.9 L1259.36 186.73 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M922.21 809.48 L894.66 809.32 L880.93 828.16 L881.74 845.78 L884.6 849.77 L922.93 857.6 L932.61 839.71 L922.21 809.48 Z"
      /><path d="M922.21 809.48 L894.66 809.32 L880.93 828.16 L881.74 845.78 L884.6 849.77 L922.93 857.6 L932.61 839.71 L922.21 809.48 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1334.5601 639.57 L1313.95 648.22 L1310.23 661.36 L1329.26 689.46 L1372.29 677.95 L1370.24 666.27 L1334.5601 639.57 Z"
      /><path d="M1334.5601 639.57 L1313.95 648.22 L1310.23 661.36 L1329.26 689.46 L1372.29 677.95 L1370.24 666.27 L1334.5601 639.57 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M84.46 313.33 L80.09 355 L41.21 346.68 L35.12 316.65 L47.72 304.12 L84.46 313.33 Z"
      /><path d="M84.46 313.33 L80.09 355 L41.21 346.68 L35.12 316.65 L47.72 304.12 L84.46 313.33 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1742.84 378.24 L1680.42 390 L1678.85 393.4 L1705.85 432.99 L1737.37 425.31 L1747.1 385.24 L1742.84 378.24 Z"
      /><path d="M1742.84 378.24 L1680.42 390 L1678.85 393.4 L1705.85 432.99 L1737.37 425.31 L1747.1 385.24 L1742.84 378.24 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M61.35 546.95 L51.32 547.29 L38.41 559.12 L37.53 573.98 L54.32 589.83 L79.98 581.27 L84 564.03 L61.35 546.95 Z"
      /><path d="M61.35 546.95 L51.32 547.29 L38.41 559.12 L37.53 573.98 L54.32 589.83 L79.98 581.27 L84 564.03 L61.35 546.95 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M867.53 127.88 L886.75 162.05 L864.47 182.76 L829.87 167.12 L829.16 165.32 L833.67 142.6 L867.53 127.88 Z"
      /><path d="M867.53 127.88 L886.75 162.05 L864.47 182.76 L829.87 167.12 L829.16 165.32 L833.67 142.6 L867.53 127.88 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M974.76 366.47 L1019.57 383.9 L996.72 430.99 L968.58 421.44 L959.35 386.96 L974.76 366.47 Z"
      /><path d="M974.76 366.47 L1019.57 383.9 L996.72 430.99 L968.58 421.44 L959.35 386.96 L974.76 366.47 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1419.4399 325.79 L1430.17 326.46 L1443.3199 370.82 L1398.83 382.64 L1393.1 345.75 L1419.4399 325.79 Z"
      /><path d="M1419.4399 325.79 L1430.17 326.46 L1443.3199 370.82 L1398.83 382.64 L1393.1 345.75 L1419.4399 325.79 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1877.5699 887.77 L1920 894.5 L1920 937.8 L1885.53 941.28 L1861.58 905.02 L1862.74 897.73 L1877.5699 887.77 Z"
      /><path d="M1877.5699 887.77 L1920 894.5 L1920 937.8 L1885.53 941.28 L1861.58 905.02 L1862.74 897.73 L1877.5699 887.77 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1222.41 100.04 L1226.0699 115.48 L1192.15 145.76 L1160.98 117.95 L1165.5699 97.6 L1200.3101 83.52 L1222.41 100.04 Z"
      /><path d="M1222.41 100.04 L1226.0699 115.48 L1192.15 145.76 L1160.98 117.95 L1165.5699 97.6 L1200.3101 83.52 L1222.41 100.04 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M362.5 256.05 L355.54 287.5 L346.14 290.12 L298.77 263.69 L297.73 255.08 L336.53 235.35 L362.5 256.05 Z"
      /><path d="M362.5 256.05 L355.54 287.5 L346.14 290.12 L298.77 263.69 L297.73 255.08 L336.53 235.35 L362.5 256.05 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1282.98 958.18 L1303.7 964.98 L1311.08 1001.67 L1305.46 1006.07 L1262.95 996.09 L1261.96 994.31 L1282.98 958.18 Z"
      /><path d="M1282.98 958.18 L1303.7 964.98 L1311.08 1001.67 L1305.46 1006.07 L1262.95 996.09 L1261.96 994.31 L1282.98 958.18 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M237.78 535.28 L207.19 534.83 L200.98 553.18 L216.25 569.85 L241.26 569.85 L248.3 546.83 L237.78 535.28 Z"
      /><path d="M237.78 535.28 L207.19 534.83 L200.98 553.18 L216.25 569.85 L241.26 569.85 L248.3 546.83 L237.78 535.28 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M531.89 137.62 L566.1 159.18 L566.1 175.01 L536.15 192.35 L516.66 170.99 L531.89 137.62 Z"
      /><path d="M531.89 137.62 L566.1 159.18 L566.1 175.01 L536.15 192.35 L516.66 170.99 L531.89 137.62 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1669.61 455.92 L1658.86 496.74 L1631.4301 490.69 L1621.99 476.46 L1629.22 450.47 L1649.01 439 L1669.61 455.92 Z"
      /><path d="M1669.61 455.92 L1658.86 496.74 L1631.4301 490.69 L1621.99 476.46 L1629.22 450.47 L1649.01 439 L1669.61 455.92 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M684.8 881.69 L644.71 890.79 L649.86 919.29 L684.44 928.07 L698.88 908.65 L684.8 881.69 Z"
      /><path d="M684.8 881.69 L644.71 890.79 L649.86 919.29 L684.44 928.07 L698.88 908.65 L684.8 881.69 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1170.8 0 L1228.9 0 L1228.26 37.17 L1200.78 52.4 L1173.0699 35.97 L1170.8 0 Z"
      /><path d="M1170.8 0 L1228.9 0 L1228.26 37.17 L1200.78 52.4 L1173.0699 35.97 L1170.8 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1204.87 659.79 L1223.02 660.41 L1246.33 684.2 L1239.04 704.5 L1214.1 706.66 L1197.38 673.94 L1204.87 659.79 Z"
      /><path d="M1204.87 659.79 L1223.02 660.41 L1246.33 684.2 L1239.04 704.5 L1214.1 706.66 L1197.38 673.94 L1204.87 659.79 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1316.11 206.44 L1284.3101 227.04 L1283.09 243.14 L1307.26 269.82 L1315.33 271.52 L1325.02 265.41 L1339.49 224.66 L1329.35 209.65 L1316.11 206.44 Z"
      /><path d="M1316.11 206.44 L1284.3101 227.04 L1283.09 243.14 L1307.26 269.82 L1315.33 271.52 L1325.02 265.41 L1339.49 224.66 L1329.35 209.65 L1316.11 206.44 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M895.3 0 L956.5 0 L956.71 10.66 L925 49.55 L903.14 44.85 L892.55 25.16 L895.3 0 Z"
      /><path d="M895.3 0 L956.5 0 L956.71 10.66 L925 49.55 L903.14 44.85 L892.55 25.16 L895.3 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M904.8 924.39 L881.11 913.5 L857.45 938.57 L864.75 950.28 L902.53 961.55 L910.29 949.36 L904.8 924.39 Z"
      /><path d="M904.8 924.39 L881.11 913.5 L857.45 938.57 L864.75 950.28 L902.53 961.55 L910.29 949.36 L904.8 924.39 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1492.2 0 L1432.1 0 L1432.09 0.23 L1455.37 59.71 L1482.29 56.07 L1496.8 33.13 L1492.2 0 Z"
      /><path d="M1492.2 0 L1432.1 0 L1432.09 0.23 L1455.37 59.71 L1482.29 56.07 L1496.8 33.13 L1492.2 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M262.99 589.74 L249.23 583.1 L216.99 614.51 L219.42 626.68 L228.11 632.16 L267.22 620.04 L262.99 589.74 Z"
      /><path d="M262.99 589.74 L249.23 583.1 L216.99 614.51 L219.42 626.68 L228.11 632.16 L267.22 620.04 L262.99 589.74 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1004.55 613.8 L1003.36 623.23 L981.35 644.98 L949.89 634.62 L938.81 598.18 L947.93 587.73 L984.45 585.74 L1004.55 613.8 Z"
      /><path d="M1004.55 613.8 L1003.36 623.23 L981.35 644.98 L949.89 634.62 L938.81 598.18 L947.93 587.73 L984.45 585.74 L1004.55 613.8 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M677.49 415.18 L657.75 428.66 L673.34 470.67 L709.51 457.91 L709.1 432.51 L677.49 415.18 Z"
      /><path d="M677.49 415.18 L657.75 428.66 L673.34 470.67 L709.51 457.91 L709.1 432.51 L677.49 415.18 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1838.7 0 L1839.22 8.9 L1809.65 43.62 L1773.5601 18.05 L1771.3 0 L1838.7 0 Z"
      /><path d="M1838.7 0 L1839.22 8.9 L1809.65 43.62 L1773.5601 18.05 L1771.3 0 L1838.7 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M560.9 0 L522.1 0 L517.93 37.77 L527.47 47.56 L562.5 33.46 L560.9 0 Z"
      /><path d="M560.9 0 L522.1 0 L517.93 37.77 L527.47 47.56 L562.5 33.46 L560.9 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M133.46 81.79 L90.17 75.96 L85.82 81.08 L97.74 131.52 L137.25 120.36 L133.46 81.79 Z"
      /><path d="M133.46 81.79 L90.17 75.96 L85.82 81.08 L97.74 131.52 L137.25 120.36 L133.46 81.79 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M19.11 370.74 L0 370.1 L0 431.9 L26.73 429.83 L37.52 390.99 L19.11 370.74 Z"
      /><path d="M19.11 370.74 L0 370.1 L0 431.9 L26.73 429.83 L37.52 390.99 L19.11 370.74 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1640.74 344.49 L1635.22 346.48 L1617.1801 380.46 L1620.84 386.35 L1675.8 394.9 L1678.85 393.4 L1680.42 390 L1676.96 366.67 L1640.74 344.49 Z"
      /><path d="M1640.74 344.49 L1635.22 346.48 L1617.1801 380.46 L1620.84 386.35 L1675.8 394.9 L1678.85 393.4 L1680.42 390 L1676.96 366.67 L1640.74 344.49 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M482.74 1017.07 L507.63 1037.78 L507.3 1080 L438.3 1080 L438.25 1041.03 L482.74 1017.07 Z"
      /><path d="M482.74 1017.07 L507.63 1037.78 L507.3 1080 L438.3 1080 L438.25 1041.03 L482.74 1017.07 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1272.05 674.12 L1278.47 676.99 L1285.9301 702.16 L1269.4 725.03 L1255.1801 726.95 L1239.04 704.5 L1246.33 684.2 L1272.05 674.12 Z"
      /><path d="M1272.05 674.12 L1278.47 676.99 L1285.9301 702.16 L1269.4 725.03 L1255.1801 726.95 L1239.04 704.5 L1246.33 684.2 L1272.05 674.12 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1741.4 567.52 L1721.12 559.36 L1683.11 564.44 L1682.01 565.16 L1674.3199 592.24 L1704.73 628.04 L1729.78 626.92 L1746.54 602.05 L1741.4 567.52 Z"
      /><path d="M1741.4 567.52 L1721.12 559.36 L1683.11 564.44 L1682.01 565.16 L1674.3199 592.24 L1704.73 628.04 L1729.78 626.92 L1746.54 602.05 L1741.4 567.52 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M996.18 906.97 L980.09 897.33 L962.43 899.65 L968.14 934.33 L983.47 939.39 L1000.13 920.84 L996.18 906.97 Z"
      /><path d="M996.18 906.97 L980.09 897.33 L962.43 899.65 L968.14 934.33 L983.47 939.39 L1000.13 920.84 L996.18 906.97 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1661.99 914.45 L1691.83 929.7 L1694.4 951.34 L1677.02 971.5 L1649.6899 968.19 L1631.3101 941.89 L1631.9301 936.44 L1661.99 914.45 Z"
      /><path d="M1661.99 914.45 L1691.83 929.7 L1694.4 951.34 L1677.02 971.5 L1649.6899 968.19 L1631.3101 941.89 L1631.9301 936.44 L1661.99 914.45 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M367.9 0 L407.8 0 L403.41 58.07 L379.28 61.24 L360.15 35.1 L367.9 0 Z"
      /><path d="M367.9 0 L407.8 0 L403.41 58.07 L379.28 61.24 L360.15 35.1 L367.9 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M228.11 632.16 L240.03 670.7 L210.79 687.05 L198.87 684.07 L184.66 647.07 L219.42 626.68 L228.11 632.16 Z"
      /><path d="M228.11 632.16 L240.03 670.7 L210.79 687.05 L198.87 684.07 L184.66 647.07 L219.42 626.68 L228.11 632.16 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M393.6 673.26 L356.94 648.7 L343.81 691.25 L359.3 702.33 L393.6 673.26 Z"
      /><path d="M393.6 673.26 L356.94 648.7 L343.81 691.25 L359.3 702.33 L393.6 673.26 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M679.61 72.31 L696.63 87.05 L685.56 125.49 L647.77 120.49 L647.01 119.64 L644.65 89.57 L679.61 72.31 Z"
      /><path d="M679.61 72.31 L696.63 87.05 L685.56 125.49 L647.77 120.49 L647.01 119.64 L644.65 89.57 L679.61 72.31 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1586.1 472.56 L1559.33 468.3 L1543.28 503.15 L1562.9399 523.64 L1585.85 512.55 L1587.24 473.81 L1586.1 472.56 Z"
      /><path d="M1586.1 472.56 L1559.33 468.3 L1543.28 503.15 L1562.9399 523.64 L1585.85 512.55 L1587.24 473.81 L1586.1 472.56 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M967.55 245.97 L952.17 241.84 L917.95 274.61 L944.58 302.65 L972.22 297.47 L981.05 283.61 L967.55 245.97 Z"
      /><path d="M967.55 245.97 L952.17 241.84 L917.95 274.61 L944.58 302.65 L972.22 297.47 L981.05 283.61 L967.55 245.97 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1821.16 109.76 L1849.27 127.73 L1840.87 166.19 L1802.0699 170.98 L1798.15 120.87 L1807.24 111.73 L1821.16 109.76 Z"
      /><path d="M1821.16 109.76 L1849.27 127.73 L1840.87 166.19 L1802.0699 170.98 L1798.15 120.87 L1807.24 111.73 L1821.16 109.76 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1689.72 866.49 L1699.75 868.54 L1718.8 904.56 L1691.83 929.7 L1661.99 914.45 L1658.83 884.39 L1689.72 866.49 Z"
      /><path d="M1689.72 866.49 L1699.75 868.54 L1718.8 904.56 L1691.83 929.7 L1661.99 914.45 L1658.83 884.39 L1689.72 866.49 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1349.42 988.6 L1381 995.82 L1373.8 1035.29 L1346.4301 1038.15 L1333.67 1003.58 L1349.42 988.6 Z"
      /><path d="M1349.42 988.6 L1381 995.82 L1373.8 1035.29 L1346.4301 1038.15 L1333.67 1003.58 L1349.42 988.6 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1788.9399 1026.83 L1824.39 1044.76 L1826.1 1080 L1769.3 1080 L1770.08 1043.25 L1788.9399 1026.83 Z"
      /><path d="M1788.9399 1026.83 L1824.39 1044.76 L1826.1 1080 L1769.3 1080 L1770.08 1043.25 L1788.9399 1026.83 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M877.51 649.41 L845.64 618.62 L824.03 628.74 L818.62 653.73 L840.07 679.27 L859.29 680.55 L877.51 649.41 Z"
      /><path d="M877.51 649.41 L845.64 618.62 L824.03 628.74 L818.62 653.73 L840.07 679.27 L859.29 680.55 L877.51 649.41 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1543.2 449.96 L1547.35 451.51 L1559.33 468.3 L1543.28 503.15 L1521.04 501.48 L1509.12 471.17 L1543.2 449.96 Z"
      /><path d="M1543.2 449.96 L1547.35 451.51 L1559.33 468.3 L1543.28 503.15 L1521.04 501.48 L1509.12 471.17 L1543.2 449.96 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1569.71 597.76 L1555.04 597.2 L1532.5699 616.7 L1533.77 641.08 L1542.27 649.24 L1584.08 647.84 L1587.48 645.32 L1590.83 626.53 L1569.71 597.76 Z"
      /><path d="M1569.71 597.76 L1555.04 597.2 L1532.5699 616.7 L1533.77 641.08 L1542.27 649.24 L1584.08 647.84 L1587.48 645.32 L1590.83 626.53 L1569.71 597.76 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1601.25 305.47 L1569.16 282.21 L1546.6801 316.56 L1578.22 340.14 L1599.84 322.16 L1601.25 305.47 Z"
      /><path d="M1601.25 305.47 L1569.16 282.21 L1546.6801 316.56 L1578.22 340.14 L1599.84 322.16 L1601.25 305.47 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1587.24 473.81 L1621.99 476.46 L1631.4301 490.69 L1607.67 519.21 L1585.85 512.55 L1587.24 473.81 Z"
      /><path d="M1587.24 473.81 L1621.99 476.46 L1631.4301 490.69 L1607.67 519.21 L1585.85 512.55 L1587.24 473.81 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M314.55 193.93 L340.18 205.31 L336.53 235.35 L297.73 255.08 L294.69 252.09 L290.01 203.54 L314.55 193.93 Z"
      /><path d="M314.55 193.93 L340.18 205.31 L336.53 235.35 L297.73 255.08 L294.69 252.09 L290.01 203.54 L314.55 193.93 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1284.3101 227.04 L1283.09 243.14 L1244.5 259.9 L1230.21 248.09 L1230.11 220.28 L1257.5699 201.83 L1284.3101 227.04 Z"
      /><path d="M1284.3101 227.04 L1283.09 243.14 L1244.5 259.9 L1230.21 248.09 L1230.11 220.28 L1257.5699 201.83 L1284.3101 227.04 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M993.19 862.59 L980.09 897.33 L962.43 899.65 L960.68 898.79 L953.81 877.1 L974.68 852.69 L993.19 862.59 Z"
      /><path d="M993.19 862.59 L980.09 897.33 L962.43 899.65 L960.68 898.79 L953.81 877.1 L974.68 852.69 L993.19 862.59 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M567.66 384.49 L594.81 403.07 L591.61 424.59 L553.73 436.71 L545.98 407.82 L567.66 384.49 Z"
      /><path d="M567.66 384.49 L594.81 403.07 L591.61 424.59 L553.73 436.71 L545.98 407.82 L567.66 384.49 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1356.74 452.47 L1343.2 443.54 L1307.8199 451.9 L1300.75 462.61 L1308.88 494.76 L1338.6 510.38 L1341.6801 508.91 L1356.74 452.47 Z"
      /><path d="M1356.74 452.47 L1343.2 443.54 L1307.8199 451.9 L1300.75 462.61 L1308.88 494.76 L1338.6 510.38 L1341.6801 508.91 L1356.74 452.47 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M309.2 0 L258.1 0 L256.9 41.73 L274.97 56.33 L315.16 43.76 L309.2 0 Z"
      /><path d="M309.2 0 L258.1 0 L256.9 41.73 L274.97 56.33 L315.16 43.76 L309.2 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M606.03 443.03 L576.22 474.94 L587.43 489.04 L628.91 476.75 L620.51 446.85 L606.03 443.03 Z"
      /><path d="M606.03 443.03 L576.22 474.94 L587.43 489.04 L628.91 476.75 L620.51 446.85 L606.03 443.03 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1214.1 706.66 L1197.38 673.94 L1170.48 685.41 L1168.42 712.26 L1189.37 729.57 L1198.74 729.21 L1214.1 706.66 Z"
      /><path d="M1214.1 706.66 L1197.38 673.94 L1170.48 685.41 L1168.42 712.26 L1189.37 729.57 L1198.74 729.21 L1214.1 706.66 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1785.01 718.38 L1812.29 724.29 L1827.27 761.98 L1799.89 789.56 L1756.61 772.72 L1764.83 729.7 L1785.01 718.38 Z"
      /><path d="M1785.01 718.38 L1812.29 724.29 L1827.27 761.98 L1799.89 789.56 L1756.61 772.72 L1764.83 729.7 L1785.01 718.38 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M960.68 898.79 L962.43 899.65 L968.14 934.33 L945.05 944.77 L943.35 943.88 L934.54 910.42 L960.68 898.79 Z"
      /><path d="M960.68 898.79 L962.43 899.65 L968.14 934.33 L945.05 944.77 L943.35 943.88 L934.54 910.42 L960.68 898.79 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1657.64 42.17 L1681.79 52.45 L1685.75 91.93 L1660.9301 101.88 L1624.17 70.68 L1657.64 42.17 Z"
      /><path d="M1657.64 42.17 L1681.79 52.45 L1685.75 91.93 L1660.9301 101.88 L1624.17 70.68 L1657.64 42.17 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1331.92 154.05 L1305.84 156.58 L1299.5 175.74 L1316.11 206.44 L1329.35 209.65 L1353.24 175.79 L1331.92 154.05 Z"
      /><path d="M1331.92 154.05 L1305.84 156.58 L1299.5 175.74 L1316.11 206.44 L1329.35 209.65 L1353.24 175.79 L1331.92 154.05 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1547.01 774.53 L1531.23 751.05 L1498.38 760.99 L1490.79 779.05 L1498.96 797.5 L1536.91 803.11 L1547.01 774.53 Z"
      /><path d="M1547.01 774.53 L1531.23 751.05 L1498.38 760.99 L1490.79 779.05 L1498.96 797.5 L1536.91 803.11 L1547.01 774.53 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M925.65 907.48 L904.8 924.39 L881.11 913.5 L879.52 890.79 L916.75 886.74 L925.65 907.48 Z"
      /><path d="M925.65 907.48 L904.8 924.39 L881.11 913.5 L879.52 890.79 L916.75 886.74 L925.65 907.48 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M730.06 908.77 L698.88 908.65 L684.44 928.07 L688.12 950.21 L731.17 960.2 L742.53 939.37 L730.06 908.77 Z"
      /><path d="M730.06 908.77 L698.88 908.65 L684.44 928.07 L688.12 950.21 L731.17 960.2 L742.53 939.37 L730.06 908.77 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M522.86 790.57 L559.85 801.51 L557.72 850.34 L551.47 854.31 L513.68 839.55 L522.86 790.57 Z"
      /><path d="M522.86 790.57 L559.85 801.51 L557.72 850.34 L551.47 854.31 L513.68 839.55 L522.86 790.57 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1019.48 885.18 L1041.4 893.66 L1041.86 895.96 L1020.96 927.31 L1000.13 920.84 L996.18 906.97 L1019.48 885.18 Z"
      /><path d="M1019.48 885.18 L1041.4 893.66 L1041.86 895.96 L1020.96 927.31 L1000.13 920.84 L996.18 906.97 L1019.48 885.18 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1526.48 269.61 L1501.17 245.07 L1483.9399 250.83 L1476.26 287.07 L1513.58 300.32 L1526.48 269.61 Z"
      /><path d="M1526.48 269.61 L1501.17 245.07 L1483.9399 250.83 L1476.26 287.07 L1513.58 300.32 L1526.48 269.61 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M483.88 695.82 L451.38 650.76 L416.9 663.88 L411.32 673.16 L415.93 690.01 L440.55 713.32 L468.08 714.33 L483.85 696.09 L483.88 695.82 Z"
      /><path d="M483.88 695.82 L451.38 650.76 L416.9 663.88 L411.32 673.16 L415.93 690.01 L440.55 713.32 L468.08 714.33 L483.85 696.09 L483.88 695.82 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1102.59 774.56 L1111.4301 775.43 L1136.13 809.13 L1102.12 833.08 L1077.47 818.44 L1074.79 807.8 L1102.59 774.56 Z"
      /><path d="M1102.59 774.56 L1111.4301 775.43 L1136.13 809.13 L1102.12 833.08 L1077.47 818.44 L1074.79 807.8 L1102.59 774.56 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1427.52 482.81 L1396.9399 505.85 L1432.27 537.64 L1443.35 534.39 L1459.6801 498.15 L1427.52 482.81 Z"
      /><path d="M1427.52 482.81 L1396.9399 505.85 L1432.27 537.64 L1443.35 534.39 L1459.6801 498.15 L1427.52 482.81 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M88.28 176.88 L80.89 211.7 L70.28 215.32 L38.77 201.36 L41.19 166.46 L42.56 165.33 L88.28 176.88 Z"
      /><path d="M88.28 176.88 L80.89 211.7 L70.28 215.32 L38.77 201.36 L41.19 166.46 L42.56 165.33 L88.28 176.88 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M983.45 762.21 L939.1 779.31 L937.97 792.54 L976.93 816.13 L988.57 809.73 L993.28 773.63 L983.45 762.21 Z"
      /><path d="M983.45 762.21 L939.1 779.31 L937.97 792.54 L976.93 816.13 L988.57 809.73 L993.28 773.63 L983.45 762.21 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M254.45 675.29 L265.77 700.95 L253.38 725.63 L225.8 733.01 L210.79 687.05 L240.03 670.7 L254.45 675.29 Z"
      /><path d="M254.45 675.29 L265.77 700.95 L253.38 725.63 L225.8 733.01 L210.79 687.05 L240.03 670.7 L254.45 675.29 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M239.96 106.08 L277.99 130.71 L278.91 151.42 L272.99 157.66 L231.25 157.86 L238.02 106.29 L239.96 106.08 Z"
      /><path d="M239.96 106.08 L277.99 130.71 L278.91 151.42 L272.99 157.66 L231.25 157.86 L238.02 106.29 L239.96 106.08 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M173.24 794.54 L141.94 817.71 L145.99 841.22 L180.3 855.2 L202.41 814.56 L193.45 801.26 L173.24 794.54 Z"
      /><path d="M173.24 794.54 L141.94 817.71 L145.99 841.22 L180.3 855.2 L202.41 814.56 L193.45 801.26 L173.24 794.54 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1659.8101 307.07 L1703.45 330.84 L1703.4399 332.07 L1676.96 366.67 L1640.74 344.49 L1659.8101 307.07 Z"
      /><path d="M1659.8101 307.07 L1703.45 330.84 L1703.4399 332.07 L1676.96 366.67 L1640.74 344.49 L1659.8101 307.07 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1045.24 1030.39 L1037.62 1037.02 L1036.1 1080 L1080.5 1080 L1082.08 1036.97 L1074.35 1030.89 L1045.24 1030.39 Z"
      /><path d="M1045.24 1030.39 L1037.62 1037.02 L1036.1 1080 L1080.5 1080 L1082.08 1036.97 L1074.35 1030.89 L1045.24 1030.39 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1002.39 1031.47 L983.58 1045.48 L984 1080 L1036.1 1080 L1037.62 1037.02 L1002.39 1031.47 Z"
      /><path d="M1002.39 1031.47 L983.58 1045.48 L984 1080 L1036.1 1080 L1037.62 1037.02 L1002.39 1031.47 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1907.3 0 L1920 0 L1920 70.5 L1894.2 56.21 L1887.22 28.46 L1907.3 0 Z"
      /><path d="M1907.3 0 L1920 0 L1920 70.5 L1894.2 56.21 L1887.22 28.46 L1907.3 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1735.46 55.24 L1711.63 36.59 L1681.79 52.45 L1685.75 91.93 L1708.21 102.79 L1713.0601 101.7 L1735.46 55.24 Z"
      /><path d="M1735.46 55.24 L1711.63 36.59 L1681.79 52.45 L1685.75 91.93 L1708.21 102.79 L1713.0601 101.7 L1735.46 55.24 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M502.95 224.37 L498.24 224.93 L494.34 229.32 L495.02 261.75 L526.08 273.91 L542.12 260.95 L540.2 247.17 L502.95 224.37 Z"
      /><path d="M502.95 224.37 L498.24 224.93 L494.34 229.32 L495.02 261.75 L526.08 273.91 L542.12 260.95 L540.2 247.17 L502.95 224.37 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M903.14 44.85 L884.22 69.05 L897.16 101.89 L914.01 105.38 L938.93 73.22 L925 49.55 L903.14 44.85 Z"
      /><path d="M903.14 44.85 L884.22 69.05 L897.16 101.89 L914.01 105.38 L938.93 73.22 L925 49.55 L903.14 44.85 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1172.9301 878.74 L1178.9301 901.87 L1158.3101 931.82 L1148.42 935.06 L1125.88 906.06 L1141.45 871.64 L1172.9301 878.74 Z"
      /><path d="M1172.9301 878.74 L1178.9301 901.87 L1158.3101 931.82 L1148.42 935.06 L1125.88 906.06 L1141.45 871.64 L1172.9301 878.74 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M522.54 560.83 L483.64 555.68 L465.9 574.22 L465.97 579.83 L498.36 605.97 L528.65 568.24 L528.58 567.54 L522.54 560.83 Z"
      /><path d="M522.54 560.83 L483.64 555.68 L465.9 574.22 L465.97 579.83 L498.36 605.97 L528.65 568.24 L528.58 567.54 L522.54 560.83 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M936.24 471.47 L912.11 485.86 L903.8 506.74 L908.74 529.58 L939.23 541.11 L972.75 524.19 L979.39 491.81 L936.24 471.47 Z"
      /><path d="M936.24 471.47 L912.11 485.86 L903.8 506.74 L908.74 529.58 L939.23 541.11 L972.75 524.19 L979.39 491.81 L936.24 471.47 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1196.86 822.41 L1183.85 830.15 L1183.26 868.8 L1225.79 870.02 L1225.73 842.92 L1196.86 822.41 Z"
      /><path d="M1196.86 822.41 L1183.85 830.15 L1183.26 868.8 L1225.79 870.02 L1225.73 842.92 L1196.86 822.41 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M680.37 164.51 L693.69 175.91 L674.46 211.8 L671.67 212.56 L659.57 209.16 L649.11 195.35 L653.69 168.06 L680.37 164.51 Z"
      /><path d="M680.37 164.51 L693.69 175.91 L674.46 211.8 L671.67 212.56 L659.57 209.16 L649.11 195.35 L653.69 168.06 L680.37 164.51 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M832.32 740.36 L816.53 728.79 L775.8 745.34 L770.76 756.84 L789.63 788.62 L825.18 781.71 L832.32 740.36 Z"
      /><path d="M832.32 740.36 L816.53 728.79 L775.8 745.34 L770.76 756.84 L789.63 788.62 L825.18 781.71 L832.32 740.36 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M272.56 299.59 L233.19 286.06 L221.27 336.96 L225.26 339.52 L267.39 337.98 L272.56 299.59 Z"
      /><path d="M272.56 299.59 L233.19 286.06 L221.27 336.96 L225.26 339.52 L267.39 337.98 L272.56 299.59 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M112.73 529.84 L125.66 538.84 L123.87 565.17 L90.45 560.05 L96.83 534.46 L112.73 529.84 Z"
      /><path d="M112.73 529.84 L125.66 538.84 L123.87 565.17 L90.45 560.05 L96.83 534.46 L112.73 529.84 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M768.1 0 L721.9 0 L720.83 33.46 L736.55 50.62 L770.4 33.42 L768.1 0 Z"
      /><path d="M768.1 0 L721.9 0 L720.83 33.46 L736.55 50.62 L770.4 33.42 L768.1 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M614.45 162.96 L606.38 186.7 L583.44 189.71 L566.1 175.01 L566.1 159.18 L594.21 134.31 L614.45 162.96 Z"
      /><path d="M614.45 162.96 L606.38 186.7 L583.44 189.71 L566.1 175.01 L566.1 159.18 L594.21 134.31 L614.45 162.96 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M554.79 359.3 L542.7 359.3 L514.05 381.91 L511.38 393.32 L513.66 398.05 L545.98 407.82 L567.66 384.49 L564.58 365.39 L554.79 359.3 Z"
      /><path d="M554.79 359.3 L542.7 359.3 L514.05 381.91 L511.38 393.32 L513.66 398.05 L545.98 407.82 L567.66 384.49 L564.58 365.39 L554.79 359.3 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1379.4301 685.07 L1372.29 677.95 L1329.26 689.46 L1320.4399 710.4 L1327.24 732.39 L1342.1 736.29 L1366.34 725.41 L1379.4399 685.11 L1379.4301 685.07 Z"
      /><path d="M1379.4301 685.07 L1372.29 677.95 L1329.26 689.46 L1320.4399 710.4 L1327.24 732.39 L1342.1 736.29 L1366.34 725.41 L1379.4399 685.11 L1379.4301 685.07 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1019.48 885.18 L1005.97 862.02 L993.19 862.59 L980.09 897.33 L996.18 906.97 L1019.48 885.18 Z"
      /><path d="M1019.48 885.18 L1005.97 862.02 L993.19 862.59 L980.09 897.33 L996.18 906.97 L1019.48 885.18 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M189.18 226.2 L223.36 269.56 L223.3 270.05 L176.21 292.73 L155.2 281.85 L151.41 246.97 L189.18 226.2 Z"
      /><path d="M189.18 226.2 L223.36 269.56 L223.3 270.05 L176.21 292.73 L155.2 281.85 L151.41 246.97 L189.18 226.2 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1030.2 946.16 L1041.51 949 L1057.75 975.91 L1038.02 994.45 L1010.54 988.64 L1007.98 964.05 L1030.2 946.16 Z"
      /><path d="M1030.2 946.16 L1041.51 949 L1057.75 975.91 L1038.02 994.45 L1010.54 988.64 L1007.98 964.05 L1030.2 946.16 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1498.28 598.89 L1486.66 601.61 L1477.99 642.06 L1489.5601 657.08 L1533.77 641.08 L1532.5699 616.7 L1498.28 598.89 Z"
      /><path d="M1498.28 598.89 L1486.66 601.61 L1477.99 642.06 L1489.5601 657.08 L1533.77 641.08 L1532.5699 616.7 L1498.28 598.89 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M402.82 573.21 L386.89 567.06 L359.64 580.4 L363.6 623.36 L398.99 621.76 L413.99 601.69 L402.82 573.21 Z"
      /><path d="M402.82 573.21 L386.89 567.06 L359.64 580.4 L363.6 623.36 L398.99 621.76 L413.99 601.69 L402.82 573.21 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M624.16 388.12 L594.81 403.07 L591.61 424.59 L606.03 443.03 L620.51 446.85 L645.17 426.9 L624.16 388.12 Z"
      /><path d="M624.16 388.12 L594.81 403.07 L591.61 424.59 L606.03 443.03 L620.51 446.85 L645.17 426.9 L624.16 388.12 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1307.26 269.82 L1283.09 243.14 L1244.5 259.9 L1247.26 284.42 L1269.62 298.37 L1307.26 269.82 Z"
      /><path d="M1307.26 269.82 L1283.09 243.14 L1244.5 259.9 L1247.26 284.42 L1269.62 298.37 L1307.26 269.82 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M650.15 961.81 L634.69 937.7 L611.45 939.11 L609.15 941.82 L615.81 984.44 L633.99 989.74 L635.2 989.26 L650.15 961.81 Z"
      /><path d="M650.15 961.81 L634.69 937.7 L611.45 939.11 L609.15 941.82 L615.81 984.44 L633.99 989.74 L635.2 989.26 L650.15 961.81 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1140.51 328.02 L1140.3101 328.1 L1128.03 344.74 L1147.9301 382.35 L1166.71 383.8 L1187.77 356.58 L1186.42 346.77 L1175.36 334.49 L1140.51 328.02 Z"
      /><path d="M1140.51 328.02 L1140.3101 328.1 L1128.03 344.74 L1147.9301 382.35 L1166.71 383.8 L1187.77 356.58 L1186.42 346.77 L1175.36 334.49 L1140.51 328.02 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M653.06 533.78 L625.07 549.59 L622.9 572.93 L626.12 578.99 L654.51 577.36 L671.28 558.67 L670.14 550.3 L653.06 533.78 Z"
      /><path d="M653.06 533.78 L625.07 549.59 L622.9 572.93 L626.12 578.99 L654.51 577.36 L671.28 558.67 L670.14 550.3 L653.06 533.78 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M918.25 383.69 L913.56 420.96 L938.12 440.17 L968.58 421.44 L959.35 386.96 L918.25 383.69 Z"
      /><path d="M918.25 383.69 L913.56 420.96 L938.12 440.17 L968.58 421.44 L959.35 386.96 L918.25 383.69 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M686.77 127.14 L680.37 164.51 L693.69 175.91 L702.6 176.55 L721.54 155.66 L717.84 134.97 L686.77 127.14 Z"
      /><path d="M686.77 127.14 L680.37 164.51 L693.69 175.91 L702.6 176.55 L721.54 155.66 L717.84 134.97 L686.77 127.14 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1255.01 820.63 L1241.62 798.67 L1201.51 807.14 L1196.86 822.41 L1225.73 842.92 L1255.01 820.63 Z"
      /><path d="M1255.01 820.63 L1241.62 798.67 L1201.51 807.14 L1196.86 822.41 L1225.73 842.92 L1255.01 820.63 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1748.97 660.26 L1779.63 665.45 L1785.01 718.38 L1764.83 729.7 L1721.49 704.34 L1721.23 700.74 L1748.97 660.26 Z"
      /><path d="M1748.97 660.26 L1779.63 665.45 L1785.01 718.38 L1764.83 729.7 L1721.49 704.34 L1721.23 700.74 L1748.97 660.26 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M588.98 351.69 L623.43 366.86 L627.61 378.97 L624.16 388.12 L594.81 403.07 L567.66 384.49 L564.58 365.39 L588.98 351.69 Z"
      /><path d="M588.98 351.69 L623.43 366.86 L627.61 378.97 L624.16 388.12 L594.81 403.07 L567.66 384.49 L564.58 365.39 L588.98 351.69 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1610.7 0 L1648.9 0 L1657.64 42.17 L1624.17 70.68 L1614.66 71.38 L1604.86 65.37 L1598.03 52.39 L1610.7 0 Z"
      /><path d="M1610.7 0 L1648.9 0 L1657.64 42.17 L1624.17 70.68 L1614.66 71.38 L1604.86 65.37 L1598.03 52.39 L1610.7 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1628.54 831.63 L1615.3101 837.22 L1599.76 874.16 L1609 888.68 L1649 879.35 L1635.51 834.15 L1628.54 831.63 Z"
      /><path d="M1628.54 831.63 L1615.3101 837.22 L1599.76 874.16 L1609 888.68 L1649 879.35 L1635.51 834.15 L1628.54 831.63 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1464.26 992.39 L1424.26 970.19 L1402.8 980.37 L1400.78 984.7 L1424.1 1028.36 L1447.71 1032.67 L1461.7 1021.32 L1464.26 992.39 Z"
      /><path d="M1464.26 992.39 L1424.26 970.19 L1402.8 980.37 L1400.78 984.7 L1424.1 1028.36 L1447.71 1032.67 L1461.7 1021.32 L1464.26 992.39 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1244.5 259.9 L1247.26 284.42 L1220.04 304.43 L1191.83 290.07 L1196.38 259.35 L1230.21 248.09 L1244.5 259.9 Z"
      /><path d="M1244.5 259.9 L1247.26 284.42 L1220.04 304.43 L1191.83 290.07 L1196.38 259.35 L1230.21 248.09 L1244.5 259.9 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M678.31 499.37 L671.49 474.05 L632.75 480.01 L632.24 506.24 L652.42 523.5 L678.31 499.37 Z"
      /><path d="M678.31 499.37 L671.49 474.05 L632.75 480.01 L632.24 506.24 L652.42 523.5 L678.31 499.37 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1734.78 491.62 L1720.85 493.59 L1717.42 497.01 L1721.12 559.36 L1741.4 567.52 L1754.4301 557.35 L1760.46 508.52 L1734.78 491.62 Z"
      /><path d="M1734.78 491.62 L1720.85 493.59 L1717.42 497.01 L1721.12 559.36 L1741.4 567.52 L1754.4301 557.35 L1760.46 508.52 L1734.78 491.62 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M75.16 664.69 L73.37 704.49 L38.99 704.4 L34.75 699.43 L42.26 668.98 L74.11 664.15 L75.16 664.69 Z"
      /><path d="M75.16 664.69 L73.37 704.49 L38.99 704.4 L34.75 699.43 L42.26 668.98 L74.11 664.15 L75.16 664.69 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M395.06 965.07 L420.13 977.33 L418.06 1021.67 L359.46 1033.09 L357.18 990.02 L395.06 965.07 Z"
      /><path d="M395.06 965.07 L420.13 977.33 L418.06 1021.67 L359.46 1033.09 L357.18 990.02 L395.06 965.07 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1065.58 283.38 L1056.35 290.69 L1058.8101 331.92 L1059.17 332.18 L1088.38 325.73 L1097.03 295.61 L1065.58 283.38 Z"
      /><path d="M1065.58 283.38 L1056.35 290.69 L1058.8101 331.92 L1059.17 332.18 L1088.38 325.73 L1097.03 295.61 L1065.58 283.38 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1631.4301 490.69 L1607.67 519.21 L1622.1801 548.17 L1644.62 544.08 L1658.9301 496.84 L1658.86 496.74 L1631.4301 490.69 Z"
      /><path d="M1631.4301 490.69 L1607.67 519.21 L1622.1801 548.17 L1644.62 544.08 L1658.9301 496.84 L1658.86 496.74 L1631.4301 490.69 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1289.79 743.38 L1269.4 725.03 L1255.1801 726.95 L1250.1801 735.56 L1258.17 771.4 L1284.02 773.12 L1289.79 743.38 Z"
      /><path d="M1289.79 743.38 L1269.4 725.03 L1255.1801 726.95 L1250.1801 735.56 L1258.17 771.4 L1284.02 773.12 L1289.79 743.38 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1189.37 729.57 L1168.42 712.26 L1134.58 725.7 L1138.3 750.84 L1166.59 764.65 L1189.37 729.57 Z"
      /><path d="M1189.37 729.57 L1168.42 712.26 L1134.58 725.7 L1138.3 750.84 L1166.59 764.65 L1189.37 729.57 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1243.16 1038.62 L1278.6899 1071.14 L1278.8 1080 L1225 1080 L1230.4 1040.89 L1243.16 1038.62 Z"
      /><path d="M1243.16 1038.62 L1278.6899 1071.14 L1278.8 1080 L1225 1080 L1230.4 1040.89 L1243.16 1038.62 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1178.9301 901.87 L1212.9399 913.57 L1199.78 953.18 L1158.3101 931.82 L1178.9301 901.87 Z"
      /><path d="M1178.9301 901.87 L1212.9399 913.57 L1199.78 953.18 L1158.3101 931.82 L1178.9301 901.87 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M611.45 939.11 L597.36 898.92 L561.23 907.15 L556.12 931.42 L570.89 952.7 L573.21 953.46 L609.15 941.82 L611.45 939.11 Z"
      /><path d="M611.45 939.11 L597.36 898.92 L561.23 907.15 L556.12 931.42 L570.89 952.7 L573.21 953.46 L609.15 941.82 L611.45 939.11 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M750.89 180.08 L778.92 187.9 L771.31 225.5 L745.46 222.01 L740.8 191.59 L750.89 180.08 Z"
      /><path d="M750.89 180.08 L778.92 187.9 L771.31 225.5 L745.46 222.01 L740.8 191.59 L750.89 180.08 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1293.51 912.83 L1277.67 948.72 L1282.98 958.18 L1303.7 964.98 L1333.96 948.61 L1326.5601 922.09 L1293.51 912.83 Z"
      /><path d="M1293.51 912.83 L1277.67 948.72 L1282.98 958.18 L1303.7 964.98 L1333.96 948.61 L1326.5601 922.09 L1293.51 912.83 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M646.99 788.19 L593.81 762.4 L581.58 791.17 L611.19 829.03 L622.13 828.84 L647.05 797.98 L646.99 788.19 Z"
      /><path d="M646.99 788.19 L593.81 762.4 L581.58 791.17 L611.19 829.03 L622.13 828.84 L647.05 797.98 L646.99 788.19 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M809.08 71.91 L793.01 61.65 L766.51 84.35 L766.15 92.92 L775.58 103.82 L814.17 105.57 L816.09 102.58 L809.08 71.91 Z"
      /><path d="M809.08 71.91 L793.01 61.65 L766.51 84.35 L766.15 92.92 L775.58 103.82 L814.17 105.57 L816.09 102.58 L809.08 71.91 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M218.83 756.49 L254.85 786.24 L227.84 819.7 L202.41 814.56 L193.45 801.26 L218.83 756.49 Z"
      /><path d="M218.83 756.49 L254.85 786.24 L227.84 819.7 L202.41 814.56 L193.45 801.26 L218.83 756.49 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1631.3101 941.89 L1649.6899 968.19 L1629.38 1000.49 L1610.45 998.31 L1590.3199 967.53 L1631.3101 941.89 Z"
      /><path d="M1631.3101 941.89 L1649.6899 968.19 L1629.38 1000.49 L1610.45 998.31 L1590.3199 967.53 L1631.3101 941.89 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M733.39 121.2 L763.11 141.46 L746.88 165.35 L721.54 155.66 L717.84 134.97 L733.39 121.2 Z"
      /><path d="M733.39 121.2 L763.11 141.46 L746.88 165.35 L721.54 155.66 L717.84 134.97 L733.39 121.2 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1629.22 450.47 L1596.64 433.25 L1586.1 472.56 L1587.24 473.81 L1621.99 476.46 L1629.22 450.47 Z"
      /><path d="M1629.22 450.47 L1596.64 433.25 L1586.1 472.56 L1587.24 473.81 L1621.99 476.46 L1629.22 450.47 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M245.17 954.12 L224.75 984.05 L172.22 969.16 L168.96 949.4 L175.39 935 L211.35 923.47 L245.17 954.12 Z"
      /><path d="M245.17 954.12 L224.75 984.05 L172.22 969.16 L168.96 949.4 L175.39 935 L211.35 923.47 L245.17 954.12 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M418.48 107.99 L452.48 114.76 L459.41 125.18 L438.35 161.08 L416.78 159.49 L410.23 114.44 L418.48 107.99 Z"
      /><path d="M418.48 107.99 L452.48 114.76 L459.41 125.18 L438.35 161.08 L416.78 159.49 L410.23 114.44 L418.48 107.99 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M864.47 182.76 L864.67 209.5 L851.83 218.36 L819.05 213.36 L813.92 198.14 L829.87 167.12 L864.47 182.76 Z"
      /><path d="M864.47 182.76 L864.67 209.5 L851.83 218.36 L819.05 213.36 L813.92 198.14 L829.87 167.12 L864.47 182.76 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M432.29 904.38 L445.94 964.58 L420.13 977.33 L395.06 965.07 L386.65 938.23 L400.96 910.48 L432.29 904.38 Z"
      /><path d="M432.29 904.38 L445.94 964.58 L420.13 977.33 L395.06 965.07 L386.65 938.23 L400.96 910.48 L432.29 904.38 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1599.98 247.03 L1624.54 259.1 L1625.61 287.58 L1601.25 305.47 L1569.16 282.21 L1565.6899 268.2 L1599.98 247.03 Z"
      /><path d="M1599.98 247.03 L1624.54 259.1 L1625.61 287.58 L1601.25 305.47 L1569.16 282.21 L1565.6899 268.2 L1599.98 247.03 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1311.08 1001.67 L1333.67 1003.58 L1346.4301 1038.15 L1334.95 1052.67 L1297.21 1038.64 L1305.46 1006.07 L1311.08 1001.67 Z"
      /><path d="M1311.08 1001.67 L1333.67 1003.58 L1346.4301 1038.15 L1334.95 1052.67 L1297.21 1038.64 L1305.46 1006.07 L1311.08 1001.67 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M44.4 0 L101.4 0 L101.48 32.57 L89.62 45.36 L50.16 32.6 L44.4 0 Z"
      /><path d="M44.4 0 L101.4 0 L101.48 32.57 L89.62 45.36 L50.16 32.6 L44.4 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M720.96 795.79 L745.77 819.34 L745.6 836.99 L726.59 858.11 L693.22 855.86 L684.07 842.62 L684.67 826.87 L712.84 797.22 L720.96 795.79 Z"
      /><path d="M720.96 795.79 L745.77 819.34 L745.6 836.99 L726.59 858.11 L693.22 855.86 L684.07 842.62 L684.67 826.87 L712.84 797.22 L720.96 795.79 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M417.28 767.92 L441.63 778.47 L455.38 809.48 L415.5 841.26 L408.31 840.08 L384.54 799.66 L386.01 792.03 L417.28 767.92 Z"
      /><path d="M417.28 767.92 L441.63 778.47 L455.38 809.48 L415.5 841.26 L408.31 840.08 L384.54 799.66 L386.01 792.03 L417.28 767.92 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1920 1032.5 L1920 1080 L1874.4 1080 L1877.12 1039.75 L1920 1032.5 Z"
      /><path d="M1920 1032.5 L1920 1080 L1874.4 1080 L1877.12 1039.75 L1920 1032.5 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M836.76 318.2 L806.88 300.97 L784.24 319.04 L788.07 354.2 L817.05 364.42 L837.35 351.49 L836.76 318.2 Z"
      /><path d="M836.76 318.2 L806.88 300.97 L784.24 319.04 L788.07 354.2 L817.05 364.42 L837.35 351.49 L836.76 318.2 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1080.78 714.46 L1040.3101 709.93 L1028.98 725.99 L1042.42 763.01 L1082.52 750.54 L1087.5699 723.77 L1080.78 714.46 Z"
      /><path d="M1080.78 714.46 L1040.3101 709.93 L1028.98 725.99 L1042.42 763.01 L1082.52 750.54 L1087.5699 723.77 L1080.78 714.46 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1418.38 916.55 L1437.28 933.22 L1424.26 970.19 L1402.8 980.37 L1377.4399 943.06 L1385.63 920.86 L1418.38 916.55 Z"
      /><path d="M1418.38 916.55 L1437.28 933.22 L1424.26 970.19 L1402.8 980.37 L1377.4399 943.06 L1385.63 920.86 L1418.38 916.55 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M284.66 912.01 L328.45 945.09 L325.44 965.51 L295.06 983.73 L253.69 952.19 L279.61 911.81 L284.66 912.01 Z"
      /><path d="M284.66 912.01 L328.45 945.09 L325.44 965.51 L295.06 983.73 L253.69 952.19 L279.61 911.81 L284.66 912.01 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M731.17 960.2 L688.12 950.21 L678.49 962.32 L683.13 990.41 L716.65 997.86 L733.75 973.92 L731.17 960.2 Z"
      /><path d="M731.17 960.2 L688.12 950.21 L678.49 962.32 L683.13 990.41 L716.65 997.86 L733.75 973.92 L731.17 960.2 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M388.43 423.74 L418.39 439.75 L409.91 473.91 L396.73 480.86 L366.76 467.25 L364.5 444.16 L388.43 423.74 Z"
      /><path d="M388.43 423.74 L418.39 439.75 L409.91 473.91 L396.73 480.86 L366.76 467.25 L364.5 444.16 L388.43 423.74 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M945.05 944.77 L943.35 943.88 L910.29 949.36 L902.53 961.55 L905.6 976.68 L921.12 989.13 L953.77 978.73 L945.05 944.77 Z"
      /><path d="M945.05 944.77 L943.35 943.88 L910.29 949.36 L902.53 961.55 L905.6 976.68 L921.12 989.13 L953.77 978.73 L945.05 944.77 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1134.58 725.7 L1127.3199 720.01 L1087.5699 723.77 L1082.52 750.54 L1102.59 774.56 L1111.4301 775.43 L1138.3 750.84 L1134.58 725.7 Z"
      /><path d="M1134.58 725.7 L1127.3199 720.01 L1087.5699 723.77 L1082.52 750.54 L1102.59 774.56 L1111.4301 775.43 L1138.3 750.84 L1134.58 725.7 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M26.73 429.83 L0 431.9 L0 481.3 L20.62 483.83 L42.96 467.45 L39.1 438.29 L26.73 429.83 Z"
      /><path d="M26.73 429.83 L0 431.9 L0 481.3 L20.62 483.83 L42.96 467.45 L39.1 438.29 L26.73 429.83 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1112.25 72.32 L1070.41 63.91 L1058.45 102.17 L1079.65 126.4 L1108.73 120.16 L1112.25 72.32 Z"
      /><path d="M1112.25 72.32 L1070.41 63.91 L1058.45 102.17 L1079.65 126.4 L1108.73 120.16 L1112.25 72.32 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M989.82 726.69 L984.42 680.39 L931.45 690.81 L944.61 727.04 L982.78 734.49 L989.82 726.69 Z"
      /><path d="M989.82 726.69 L984.42 680.39 L931.45 690.81 L944.61 727.04 L982.78 734.49 L989.82 726.69 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M73.37 704.49 L81.73 712.01 L67.92 746.7 L37.9 731.92 L38.99 704.4 L73.37 704.49 Z"
      /><path d="M73.37 704.49 L81.73 712.01 L67.92 746.7 L37.9 731.92 L38.99 704.4 L73.37 704.49 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M320.97 323.75 L285.94 292.46 L272.56 299.59 L267.39 337.98 L271.25 342.21 L301 346.71 L320.99 324.12 L320.97 323.75 Z"
      /><path d="M320.97 323.75 L285.94 292.46 L272.56 299.59 L267.39 337.98 L271.25 342.21 L301 346.71 L320.99 324.12 L320.97 323.75 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1621.87 663.8 L1615.59 699.49 L1576.27 697.03 L1584.08 647.84 L1587.48 645.32 L1621.87 663.8 Z"
      /><path d="M1621.87 663.8 L1615.59 699.49 L1576.27 697.03 L1584.08 647.84 L1587.48 645.32 L1621.87 663.8 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M343.1 932.3 L386.65 938.23 L395.06 965.07 L357.18 990.02 L325.44 965.51 L328.45 945.09 L343.1 932.3 Z"
      /><path d="M343.1 932.3 L386.65 938.23 L395.06 965.07 L357.18 990.02 L325.44 965.51 L328.45 945.09 L343.1 932.3 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M807.17 841.91 L783.91 860.82 L780.64 887.05 L792.56 901.89 L826.23 901.28 L838.52 884.17 L835.41 859.21 L821.69 842.89 L807.17 841.91 Z"
      /><path d="M807.17 841.91 L783.91 860.82 L780.64 887.05 L792.56 901.89 L826.23 901.28 L838.52 884.17 L835.41 859.21 L821.69 842.89 L807.17 841.91 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1346.76 812.98 L1379.0601 824.62 L1375.4399 852.93 L1329.34 865.52 L1328.86 865.23 L1317.04 839.46 L1346.76 812.98 Z"
      /><path d="M1346.76 812.98 L1379.0601 824.62 L1375.4399 852.93 L1329.34 865.52 L1328.86 865.23 L1317.04 839.46 L1346.76 812.98 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1147.22 1037.3199 L1128.62 1051.97 L1127.1 1080 L1181 1080 L1179 1048.79 L1168.14 1038.9301 L1147.22 1037.3199 Z"
      /><path d="M1147.22 1037.3199 L1128.62 1051.97 L1127.1 1080 L1181 1080 L1179 1048.79 L1168.14 1038.9301 L1147.22 1037.3199 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M542.7 359.3 L514.05 381.91 L492.28 346.4 L516.77 333.37 L542.7 359.3 Z"
      /><path d="M542.7 359.3 L514.05 381.91 L492.28 346.4 L516.77 333.37 L542.7 359.3 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1093.9399 527.93 L1089.5 528.79 L1066.76 568.26 L1107.65 595.4 L1115.96 588.32 L1115.49 543.31 L1093.9399 527.93 Z"
      /><path d="M1093.9399 527.93 L1089.5 528.79 L1066.76 568.26 L1107.65 595.4 L1115.96 588.32 L1115.49 543.31 L1093.9399 527.93 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M97.36 132.02 L49.25 130.53 L42.56 165.33 L88.28 176.88 L98.49 168.81 L97.36 132.02 Z"
      /><path d="M97.36 132.02 L49.25 130.53 L42.56 165.33 L88.28 176.88 L98.49 168.81 L97.36 132.02 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1284 0 L1286.88 22.57 L1316.4 44.46 L1355 2.45 L1355 0 L1284 0 Z"
      /><path d="M1284 0 L1286.88 22.57 L1316.4 44.46 L1355 2.45 L1355 0 L1284 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M402.77 250.57 L388.62 243.38 L362.5 256.05 L355.54 287.5 L374.39 301.88 L383.11 302.43 L414.86 281.7 L402.77 250.57 Z"
      /><path d="M402.77 250.57 L388.62 243.38 L362.5 256.05 L355.54 287.5 L374.39 301.88 L383.11 302.43 L414.86 281.7 L402.77 250.57 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M411.32 673.16 L415.93 690.01 L382.83 728.75 L368.32 727.8 L359.3 702.33 L393.6 673.26 L411.32 673.16 Z"
      /><path d="M411.32 673.16 L415.93 690.01 L382.83 728.75 L368.32 727.8 L359.3 702.33 L393.6 673.26 L411.32 673.16 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M345.91 484.61 L317.71 478.3 L306.12 488.08 L301.9 507.45 L322.6 534.97 L332.53 537.24 L354.28 521.07 L345.91 484.61 Z"
      /><path d="M345.91 484.61 L317.71 478.3 L306.12 488.08 L301.9 507.45 L322.6 534.97 L332.53 537.24 L354.28 521.07 L345.91 484.61 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1446.8199 693.29 L1457.15 695.82 L1474.9 726.32 L1445.17 750.44 L1417.35 737.13 L1418.3101 716.35 L1446.8199 693.29 Z"
      /><path d="M1446.8199 693.29 L1457.15 695.82 L1474.9 726.32 L1445.17 750.44 L1417.35 737.13 L1418.3101 716.35 L1446.8199 693.29 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1677.02 971.5 L1649.6899 968.19 L1629.38 1000.49 L1640.92 1016.11 L1674.46 1015.79 L1684.95 998.44 L1677.02 971.5 Z"
      /><path d="M1677.02 971.5 L1649.6899 968.19 L1629.38 1000.49 L1640.92 1016.11 L1674.46 1015.79 L1684.95 998.44 L1677.02 971.5 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1693.27 155.34 L1685.42 157.97 L1671.1899 194.81 L1694.4301 217.74 L1734.53 209.06 L1734.89 208.17 L1721.6 164.96 L1693.27 155.34 Z"
      /><path d="M1693.27 155.34 L1685.42 157.97 L1671.1899 194.81 L1694.4301 217.74 L1734.53 209.06 L1734.89 208.17 L1721.6 164.96 L1693.27 155.34 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M497 628.24 L508.44 668.63 L483.88 695.82 L451.38 650.76 L456.22 640.31 L497 628.24 Z"
      /><path d="M497 628.24 L508.44 668.63 L483.88 695.82 L451.38 650.76 L456.22 640.31 L497 628.24 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1685.42 157.97 L1671.1899 194.81 L1643.22 201.78 L1627.9399 194.15 L1620.17 172.24 L1637.29 139.33 L1649.3199 135.7 L1685.42 157.97 Z"
      /><path d="M1685.42 157.97 L1671.1899 194.81 L1643.22 201.78 L1627.9399 194.15 L1620.17 172.24 L1637.29 139.33 L1649.3199 135.7 L1685.42 157.97 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1492.2 0 L1554 0 L1550.71 37.38 L1544.77 42.56 L1496.8 33.13 L1492.2 0 Z"
      /><path d="M1492.2 0 L1554 0 L1550.71 37.38 L1544.77 42.56 L1496.8 33.13 L1492.2 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M215.59 404.28 L192.2 387.02 L158.05 393.14 L150.27 406.01 L175.47 444.2 L216.17 408.5 L215.59 404.28 Z"
      /><path d="M215.59 404.28 L192.2 387.02 L158.05 393.14 L150.27 406.01 L175.47 444.2 L216.17 408.5 L215.59 404.28 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M314.36 157.28 L314.55 193.93 L290.01 203.54 L277.01 197.21 L272.99 157.66 L278.91 151.42 L314.36 157.28 Z"
      /><path d="M314.36 157.28 L314.55 193.93 L290.01 203.54 L277.01 197.21 L272.99 157.66 L278.91 151.42 L314.36 157.28 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1689.72 866.49 L1670.9301 823.76 L1635.51 834.15 L1649 879.35 L1658.83 884.39 L1689.72 866.49 Z"
      /><path d="M1689.72 866.49 L1670.9301 823.76 L1635.51 834.15 L1649 879.35 L1658.83 884.39 L1689.72 866.49 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1804.5601 812.33 L1783.5699 839.97 L1809.0699 876.86 L1830.8 872.28 L1846.54 830.24 L1804.5601 812.33 Z"
      /><path d="M1804.5601 812.33 L1783.5699 839.97 L1809.0699 876.86 L1830.8 872.28 L1846.54 830.24 L1804.5601 812.33 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M486.48 437.54 L461.13 408.55 L441.66 412.86 L430.58 434.5 L462.49 460.86 L482.72 447.92 L486.48 437.54 Z"
      /><path d="M486.48 437.54 L461.13 408.55 L441.66 412.86 L430.58 434.5 L462.49 460.86 L482.72 447.92 L486.48 437.54 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M622.13 828.84 L641.24 851.76 L636.49 883.97 L603.56 889.34 L587.79 853.63 L611.19 829.03 L622.13 828.84 Z"
      /><path d="M622.13 828.84 L641.24 851.76 L636.49 883.97 L603.56 889.34 L587.79 853.63 L611.19 829.03 L622.13 828.84 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M842.5 934.86 L857.45 938.57 L864.75 950.28 L851.48 1006.7 L807.29 963.98 L842.5 934.86 Z"
      /><path d="M842.5 934.86 L857.45 938.57 L864.75 950.28 L851.48 1006.7 L807.29 963.98 L842.5 934.86 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1920 287.1 L1920 226.4 L1875.01 228.34 L1870.62 287.28 L1878.89 291.32 L1920 287.1 Z"
      /><path d="M1920 287.1 L1920 226.4 L1875.01 228.34 L1870.62 287.28 L1878.89 291.32 L1920 287.1 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1658.9301 496.84 L1687.22 506.56 L1683.11 564.44 L1682.01 565.16 L1644.62 544.08 L1658.9301 496.84 Z"
      /><path d="M1658.9301 496.84 L1687.22 506.56 L1683.11 564.44 L1682.01 565.16 L1644.62 544.08 L1658.9301 496.84 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1920 937.8 L1920 994.7 L1883.04 988.7 L1871.77 962.79 L1885.53 941.28 L1920 937.8 Z"
      /><path d="M1920 937.8 L1920 994.7 L1883.04 988.7 L1871.77 962.79 L1885.53 941.28 L1920 937.8 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M669.94 254.08 L694.27 258.92 L700.68 290.37 L698.14 295.6 L655.9 294.31 L650.55 288.65 L650.41 287.31 L665.99 255.76 L669.94 254.08 Z"
      /><path d="M669.94 254.08 L694.27 258.92 L700.68 290.37 L698.14 295.6 L655.9 294.31 L650.55 288.65 L650.41 287.31 L665.99 255.76 L669.94 254.08 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M84.67 467.94 L61.76 476.13 L61.05 505.76 L77.76 515.25 L97.23 497.89 L91.3 472.64 L84.67 467.94 Z"
      /><path d="M84.67 467.94 L61.76 476.13 L61.05 505.76 L77.76 515.25 L97.23 497.89 L91.3 472.64 L84.67 467.94 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M511.38 393.32 L513.66 398.05 L503.77 428.49 L486.48 437.54 L461.13 408.55 L472.55 390.49 L511.38 393.32 Z"
      /><path d="M511.38 393.32 L513.66 398.05 L503.77 428.49 L486.48 437.54 L461.13 408.55 L472.55 390.49 L511.38 393.32 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1580.21 964.78 L1563.1801 975.38 L1557.78 1024.0601 L1564.11 1029.52 L1586.51 1028.11 L1610.45 998.31 L1590.3199 967.53 L1580.21 964.78 Z"
      /><path d="M1580.21 964.78 L1563.1801 975.38 L1557.78 1024.0601 L1564.11 1029.52 L1586.51 1028.11 L1610.45 998.31 L1590.3199 967.53 L1580.21 964.78 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M736.55 50.62 L720.83 33.46 L678.81 46.7 L679.61 72.31 L696.63 87.05 L713.58 85.72 L736.7 55.72 L736.55 50.62 Z"
      /><path d="M736.55 50.62 L720.83 33.46 L678.81 46.7 L679.61 72.31 L696.63 87.05 L713.58 85.72 L736.7 55.72 L736.55 50.62 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1799.89 789.56 L1756.61 772.72 L1754.88 773.69 L1737.1899 830.44 L1739.13 835.86 L1752.73 843.92 L1783.5699 839.97 L1804.5601 812.33 L1799.89 789.56 Z"
      /><path d="M1799.89 789.56 L1756.61 772.72 L1754.88 773.69 L1737.1899 830.44 L1739.13 835.86 L1752.73 843.92 L1783.5699 839.97 L1804.5601 812.33 L1799.89 789.56 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1223.7 488.04 L1213.23 513.76 L1197.17 517.92 L1163.72 487.98 L1171.85 469.55 L1209.3199 465.89 L1223.7 488.04 Z"
      /><path d="M1223.7 488.04 L1213.23 513.76 L1197.17 517.92 L1163.72 487.98 L1171.85 469.55 L1209.3199 465.89 L1223.7 488.04 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M588.26 504.44 L605.5 519.91 L605.73 532.69 L578.67 553.44 L565.74 546.27 L560.5 523.59 L588.26 504.44 Z"
      /><path d="M588.26 504.44 L605.5 519.91 L605.73 532.69 L578.67 553.44 L565.74 546.27 L560.5 523.59 L588.26 504.44 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1313.59 351.51 L1346.84 357.43 L1355.6801 389.41 L1340.59 403.63 L1306.09 395.11 L1299.5 369.69 L1313.59 351.51 Z"
      /><path d="M1313.59 351.51 L1346.84 357.43 L1355.6801 389.41 L1340.59 403.63 L1306.09 395.11 L1299.5 369.69 L1313.59 351.51 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1402.8 980.37 L1377.4399 943.06 L1342.6801 953.44 L1349.42 988.6 L1381 995.82 L1400.78 984.7 L1402.8 980.37 Z"
      /><path d="M1402.8 980.37 L1377.4399 943.06 L1342.6801 953.44 L1349.42 988.6 L1381 995.82 L1400.78 984.7 L1402.8 980.37 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1433.16 226.39 L1426.0699 175.24 L1384.04 187.96 L1384.1899 224 L1433.16 226.39 Z"
      /><path d="M1433.16 226.39 L1426.0699 175.24 L1384.04 187.96 L1384.1899 224 L1433.16 226.39 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1631.9301 936.44 L1605.0699 907.6 L1570.7 923.06 L1580.21 964.78 L1590.3199 967.53 L1631.3101 941.89 L1631.9301 936.44 Z"
      /><path d="M1631.9301 936.44 L1605.0699 907.6 L1570.7 923.06 L1580.21 964.78 L1590.3199 967.53 L1631.3101 941.89 L1631.9301 936.44 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M636.09 612.09 L617.88 629.23 L621.76 640.02 L658.71 648.64 L661.32 616.96 L636.09 612.09 Z"
      /><path d="M636.09 612.09 L617.88 629.23 L621.76 640.02 L658.71 648.64 L661.32 616.96 L636.09 612.09 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M636.09 612.09 L625.73 580.36 L599.07 602.77 L602.99 622.43 L617.88 629.23 L636.09 612.09 Z"
      /><path d="M636.09 612.09 L625.73 580.36 L599.07 602.77 L602.99 622.43 L617.88 629.23 L636.09 612.09 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1192.04 783.43 L1171 775.25 L1143.8 810.8 L1152.78 822.52 L1183.85 830.15 L1196.86 822.41 L1201.51 807.14 L1192.04 783.43 Z"
      /><path d="M1192.04 783.43 L1171 775.25 L1143.8 810.8 L1152.78 822.52 L1183.85 830.15 L1196.86 822.41 L1201.51 807.14 L1192.04 783.43 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M813.08 459.91 L840.16 473.4 L845.17 497.66 L835.03 518.61 L798.01 524.54 L778.44 511.21 L789.84 469.84 L813.08 459.91 Z"
      /><path d="M813.08 459.91 L840.16 473.4 L845.17 497.66 L835.03 518.61 L798.01 524.54 L778.44 511.21 L789.84 469.84 L813.08 459.91 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M396.22 168.86 L376.64 135.05 L347.28 154.79 L357.43 174.82 L396.22 168.86 Z"
      /><path d="M396.22 168.86 L376.64 135.05 L347.28 154.79 L357.43 174.82 L396.22 168.86 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M458.9 475.46 L490.43 502.02 L490.63 511.49 L480.66 522.49 L440.27 520.9 L440.49 488.16 L458.9 475.46 Z"
      /><path d="M458.9 475.46 L490.43 502.02 L490.63 511.49 L480.66 522.49 L440.27 520.9 L440.49 488.16 L458.9 475.46 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M348.85 200.54 L340.18 205.31 L336.53 235.35 L362.5 256.05 L388.62 243.38 L385.96 213.95 L348.85 200.54 Z"
      /><path d="M348.85 200.54 L340.18 205.31 L336.53 235.35 L362.5 256.05 L388.62 243.38 L385.96 213.95 L348.85 200.54 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M89.96 617.71 L104.42 636.37 L85.62 663.37 L75.16 664.69 L74.11 664.15 L63.2 625.96 L89.96 617.71 Z"
      /><path d="M89.96 617.71 L104.42 636.37 L85.62 663.37 L75.16 664.69 L74.11 664.15 L63.2 625.96 L89.96 617.71 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1907.3 0 L1838.7 0 L1839.22 8.9 L1856.4 28.65 L1887.22 28.46 L1907.3 0 Z"
      /><path d="M1907.3 0 L1838.7 0 L1839.22 8.9 L1856.4 28.65 L1887.22 28.46 L1907.3 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1870.62 287.28 L1848.23 292.33 L1837.28 337.23 L1865.73 359.89 L1887.2 345.36 L1878.89 291.32 L1870.62 287.28 Z"
      /><path d="M1870.62 287.28 L1848.23 292.33 L1837.28 337.23 L1865.73 359.89 L1887.2 345.36 L1878.89 291.32 L1870.62 287.28 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M445.94 964.58 L456.77 966.23 L483.66 994.61 L482.74 1017.07 L438.25 1041.03 L418.06 1021.67 L420.13 977.33 L445.94 964.58 Z"
      /><path d="M445.94 964.58 L456.77 966.23 L483.66 994.61 L482.74 1017.07 L438.25 1041.03 L418.06 1021.67 L420.13 977.33 L445.94 964.58 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M0 698.2 L0 744.3 L18.75 746.32 L37.9 731.92 L38.99 704.4 L34.75 699.43 L0 698.2 Z"
      /><path d="M0 698.2 L0 744.3 L18.75 746.32 L37.9 731.92 L38.99 704.4 L34.75 699.43 L0 698.2 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1018.94 822.52 L988.57 809.73 L976.93 816.13 L968.72 838.72 L974.68 852.69 L993.19 862.59 L1005.97 862.02 L1024.46 838.68 L1018.94 822.52 Z"
      /><path d="M1018.94 822.52 L988.57 809.73 L976.93 816.13 L968.72 838.72 L974.68 852.69 L993.19 862.59 L1005.97 862.02 L1024.46 838.68 L1018.94 822.52 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1586.51 1028.11 L1613.15 1052.92 L1609.1 1080 L1558.5 1080 L1564.11 1029.52 L1586.51 1028.11 Z"
      /><path d="M1586.51 1028.11 L1613.15 1052.92 L1609.1 1080 L1558.5 1080 L1564.11 1029.52 L1586.51 1028.11 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1682.91 1039.1801 L1716.08 1045.41 L1720.1 1080 L1666.2 1080 L1665.23 1063.58 L1682.91 1039.1801 Z"
      /><path d="M1682.91 1039.1801 L1716.08 1045.41 L1720.1 1080 L1666.2 1080 L1665.23 1063.58 L1682.91 1039.1801 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M121.68 302.89 L104.94 298.43 L84.46 313.33 L80.09 355 L89.08 368.52 L94.43 369.47 L136.95 347.25 L121.68 302.89 Z"
      /><path d="M121.68 302.89 L104.94 298.43 L84.46 313.33 L80.09 355 L89.08 368.52 L94.43 369.47 L136.95 347.25 L121.68 302.89 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1057.75 975.91 L1038.02 994.45 L1045.24 1030.39 L1074.35 1030.89 L1081.6801 989.5 L1070.26 977.26 L1057.75 975.91 Z"
      /><path d="M1057.75 975.91 L1038.02 994.45 L1045.24 1030.39 L1074.35 1030.89 L1081.6801 989.5 L1070.26 977.26 L1057.75 975.91 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M565.52 1046.7 L560.8 1080 L507.3 1080 L507.63 1037.78 L544.19 1022.5 L565.52 1046.7 Z"
      /><path d="M565.52 1046.7 L560.8 1080 L507.3 1080 L507.63 1037.78 L544.19 1022.5 L565.52 1046.7 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M817.05 364.42 L819.78 407.99 L812.22 414.83 L769.89 409.54 L768.9 367.18 L788.07 354.2 L817.05 364.42 Z"
      /><path d="M817.05 364.42 L819.78 407.99 L812.22 414.83 L769.89 409.54 L768.9 367.18 L788.07 354.2 L817.05 364.42 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1199.78 953.18 L1158.3101 931.82 L1148.42 935.06 L1142.79 946.05 L1165.23 987.42 L1178.4301 990.89 L1201.67 957.84 L1199.78 953.18 Z"
      /><path d="M1199.78 953.18 L1158.3101 931.82 L1148.42 935.06 L1142.79 946.05 L1165.23 987.42 L1178.4301 990.89 L1201.67 957.84 L1199.78 953.18 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1138.6801 265.9 L1124.89 262.55 L1122.62 263.84 L1106.86 291.26 L1140.3101 328.1 L1140.51 328.02 L1155.96 288.74 L1138.6801 265.9 Z"
      /><path d="M1138.6801 265.9 L1124.89 262.55 L1122.62 263.84 L1106.86 291.26 L1140.3101 328.1 L1140.51 328.02 L1155.96 288.74 L1138.6801 265.9 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M108.59 922.12 L78.39 895.87 L56.19 900.29 L44 926.65 L55.14 947.88 L105.46 946.86 L108.34 942.55 L108.59 922.12 Z"
      /><path d="M108.59 922.12 L78.39 895.87 L56.19 900.29 L44 926.65 L55.14 947.88 L105.46 946.86 L108.34 942.55 L108.59 922.12 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1764.83 729.7 L1756.61 772.72 L1754.88 773.69 L1709.9301 766.03 L1695.37 741.63 L1696.33 732.66 L1721.49 704.34 L1764.83 729.7 Z"
      /><path d="M1764.83 729.7 L1756.61 772.72 L1754.88 773.69 L1709.9301 766.03 L1695.37 741.63 L1696.33 732.66 L1721.49 704.34 L1764.83 729.7 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1102.59 1034.1899 L1128.62 1051.97 L1127.1 1080 L1080.5 1080 L1082.08 1036.97 L1102.59 1034.1899 Z"
      /><path d="M1102.59 1034.1899 L1128.62 1051.97 L1127.1 1080 L1080.5 1080 L1082.08 1036.97 L1102.59 1034.1899 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1754.88 773.69 L1737.1899 830.44 L1689.51 804.28 L1709.9301 766.03 L1754.88 773.69 Z"
      /><path d="M1754.88 773.69 L1737.1899 830.44 L1689.51 804.28 L1709.9301 766.03 L1754.88 773.69 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1887.22 28.46 L1856.4 28.65 L1853.9399 68.19 L1856.04 69.2 L1894.2 56.21 L1887.22 28.46 Z"
      /><path d="M1887.22 28.46 L1856.4 28.65 L1853.9399 68.19 L1856.04 69.2 L1894.2 56.21 L1887.22 28.46 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1228.23 965.84 L1237.03 985.87 L1213.87 1013.05 L1179.35 992.63 L1178.4301 990.89 L1201.67 957.84 L1228.23 965.84 Z"
      /><path d="M1228.23 965.84 L1237.03 985.87 L1213.87 1013.05 L1179.35 992.63 L1178.4301 990.89 L1201.67 957.84 L1228.23 965.84 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1160.48 442.07 L1126.67 433.27 L1105.99 468.44 L1115.64 488.17 L1149.9 495.53 L1163.72 487.98 L1171.85 469.55 L1160.48 442.07 Z"
      /><path d="M1160.48 442.07 L1126.67 433.27 L1105.99 468.44 L1115.64 488.17 L1149.9 495.53 L1163.72 487.98 L1171.85 469.55 L1160.48 442.07 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M949.89 634.62 L981.35 644.98 L986.05 677.94 L984.42 680.39 L931.45 690.81 L927.54 688.37 L921.71 662.31 L949.89 634.62 Z"
      /><path d="M949.89 634.62 L981.35 644.98 L986.05 677.94 L984.42 680.39 L931.45 690.81 L927.54 688.37 L921.71 662.31 L949.89 634.62 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M769.89 409.54 L812.22 414.83 L813.08 459.91 L789.84 469.84 L760.99 451.67 L758.64 418.47 L769.89 409.54 Z"
      /><path d="M769.89 409.54 L812.22 414.83 L813.08 459.91 L789.84 469.84 L760.99 451.67 L758.64 418.47 L769.89 409.54 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M386.01 792.03 L350.73 759.7 L323.42 784.99 L322.74 801.23 L342.21 821.47 L384.54 799.66 L386.01 792.03 Z"
      /><path d="M386.01 792.03 L350.73 759.7 L323.42 784.99 L322.74 801.23 L342.21 821.47 L384.54 799.66 L386.01 792.03 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M433.19 549.52 L465.9 574.22 L465.97 579.83 L442.38 605.9 L413.99 601.69 L402.82 573.21 L433.19 549.52 Z"
      /><path d="M433.19 549.52 L465.9 574.22 L465.97 579.83 L442.38 605.9 L413.99 601.69 L402.82 573.21 L433.19 549.52 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1163.71 598.67 L1160.4 631.16 L1147.47 640.99 L1102.33 619.32 L1107.65 595.4 L1115.96 588.32 L1152.26 586.65 L1163.71 598.67 Z"
      /><path d="M1163.71 598.67 L1160.4 631.16 L1147.47 640.99 L1102.33 619.32 L1107.65 595.4 L1115.96 588.32 L1152.26 586.65 L1163.71 598.67 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M277.01 197.21 L290.01 203.54 L294.69 252.09 L248.71 245.48 L245.73 207.9 L277.01 197.21 Z"
      /><path d="M277.01 197.21 L290.01 203.54 L294.69 252.09 L248.71 245.48 L245.73 207.9 L277.01 197.21 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1476.26 287.07 L1513.58 300.32 L1521.74 319.76 L1482.8 338.56 L1452.89 310.4 L1455.78 299.92 L1476.26 287.07 Z"
      /><path d="M1476.26 287.07 L1513.58 300.32 L1521.74 319.76 L1482.8 338.56 L1452.89 310.4 L1455.78 299.92 L1476.26 287.07 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M149.79 661.02 L155.57 693.74 L128.51 698.36 L112.05 684.53 L111.16 679.68 L133.73 655.33 L149.79 661.02 Z"
      /><path d="M149.79 661.02 L155.57 693.74 L128.51 698.36 L112.05 684.53 L111.16 679.68 L133.73 655.33 L149.79 661.02 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M996.72 430.99 L1001.96 440.1 L988.24 486.52 L979.39 491.81 L936.24 471.47 L938.12 440.17 L968.58 421.44 L996.72 430.99 Z"
      /><path d="M996.72 430.99 L1001.96 440.1 L988.24 486.52 L979.39 491.81 L936.24 471.47 L938.12 440.17 L968.58 421.44 L996.72 430.99 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M881.74 845.78 L884.6 849.77 L879.04 890.19 L838.52 884.17 L835.41 859.21 L881.74 845.78 Z"
      /><path d="M881.74 845.78 L884.6 849.77 L879.04 890.19 L838.52 884.17 L835.41 859.21 L881.74 845.78 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1607.83 117.67 L1575.74 129.81 L1580.85 163.09 L1620.17 172.24 L1637.29 139.33 L1607.83 117.67 Z"
      /><path d="M1607.83 117.67 L1575.74 129.81 L1580.85 163.09 L1620.17 172.24 L1637.29 139.33 L1607.83 117.67 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1385.4301 280.58 L1383.7 280.18 L1359.61 316.26 L1364.64 335.87 L1393.1 345.75 L1419.4399 325.79 L1385.4301 280.58 Z"
      /><path d="M1385.4301 280.58 L1383.7 280.18 L1359.61 316.26 L1364.64 335.87 L1393.1 345.75 L1419.4399 325.79 L1385.4301 280.58 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M377.79 862.57 L374.42 881.95 L345.01 895.39 L323.48 883.01 L318.17 858.37 L341.86 836.34 L377.79 862.57 Z"
      /><path d="M377.79 862.57 L374.42 881.95 L345.01 895.39 L323.48 883.01 L318.17 858.37 L341.86 836.34 L377.79 862.57 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M938.93 73.22 L966.81 77.92 L975.02 89.76 L959.39 135.15 L957 136.4 L930.18 131.54 L914.01 105.38 L938.93 73.22 Z"
      /><path d="M938.93 73.22 L966.81 77.92 L975.02 89.76 L959.39 135.15 L957 136.4 L930.18 131.54 L914.01 105.38 L938.93 73.22 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1274.03 318.52 L1308.17 327.93 L1313.59 351.51 L1299.5 369.69 L1270.79 364.93 L1257.58 339.88 L1274.03 318.52 Z"
      /><path d="M1274.03 318.52 L1308.17 327.93 L1313.59 351.51 L1299.5 369.69 L1270.79 364.93 L1257.58 339.88 L1274.03 318.52 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1480.24 362.57 L1515.95 374.92 L1517.8 387.69 L1494.58 416.59 L1459.28 381.03 L1459.1899 380.18 L1480.24 362.57 Z"
      /><path d="M1480.24 362.57 L1515.95 374.92 L1517.8 387.69 L1494.58 416.59 L1459.28 381.03 L1459.1899 380.18 L1480.24 362.57 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M143.75 349.94 L136.95 347.25 L94.43 369.47 L123.88 412.87 L150.27 406.01 L158.05 393.14 L143.75 349.94 Z"
      /><path d="M143.75 349.94 L136.95 347.25 L94.43 369.47 L123.88 412.87 L150.27 406.01 L158.05 393.14 L143.75 349.94 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1023.43 288.52 L1016.47 280.2 L981.05 283.61 L972.22 297.47 L989.9 329.61 L1018.03 328.21 L1023.43 288.52 Z"
      /><path d="M1023.43 288.52 L1016.47 280.2 L981.05 283.61 L972.22 297.47 L989.9 329.61 L1018.03 328.21 L1023.43 288.52 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1756.09 895.2 L1795.61 898.36 L1806.26 928.94 L1783.37 949.91 L1752.3199 943.73 L1741.7 907.94 L1756.09 895.2 Z"
      /><path d="M1756.09 895.2 L1795.61 898.36 L1806.26 928.94 L1783.37 949.91 L1752.3199 943.73 L1741.7 907.94 L1756.09 895.2 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M784.24 319.04 L755.29 308.93 L733.03 329.54 L731.27 352.79 L733.23 356.72 L768.9 367.18 L788.07 354.2 L784.24 319.04 Z"
      /><path d="M784.24 319.04 L755.29 308.93 L733.03 329.54 L731.27 352.79 L733.23 356.72 L768.9 367.18 L788.07 354.2 L784.24 319.04 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M316.26 44.51 L315.16 43.76 L274.97 56.33 L274.35 79.86 L301.85 103.1 L323.82 89.61 L328.15 78.14 L316.26 44.51 Z"
      /><path d="M316.26 44.51 L315.16 43.76 L274.97 56.33 L274.35 79.86 L301.85 103.1 L323.82 89.61 L328.15 78.14 L316.26 44.51 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M776.45 995.01 L733.75 973.92 L716.65 997.86 L720.88 1024.34 L731.27 1031.6801 L769.07 1026.8101 L778.2 1016.46 L776.45 995.01 Z"
      /><path d="M776.45 995.01 L733.75 973.92 L716.65 997.86 L720.88 1024.34 L731.27 1031.6801 L769.07 1026.8101 L778.2 1016.46 L776.45 995.01 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1285.26 93.47 L1303.9301 110.89 L1297.61 144.82 L1254.64 141.09 L1249.65 129.63 L1285.26 93.47 Z"
      /><path d="M1285.26 93.47 L1303.9301 110.89 L1297.61 144.82 L1254.64 141.09 L1249.65 129.63 L1285.26 93.47 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M37.53 573.98 L0 593.4 L0 602.6 L43.3 622.13 L49.47 619.61 L54.32 589.83 L37.53 573.98 Z"
      /><path d="M37.53 573.98 L0 593.4 L0 602.6 L43.3 622.13 L49.47 619.61 L54.32 589.83 L37.53 573.98 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M263.72 465.47 L231.32 452.54 L217.26 464.71 L214.8 486.24 L221.03 494.45 L244.34 502.07 L253.38 498.8 L265.48 471.98 L263.72 465.47 Z"
      /><path d="M263.72 465.47 L231.32 452.54 L217.26 464.71 L214.8 486.24 L221.03 494.45 L244.34 502.07 L253.38 498.8 L265.48 471.98 L263.72 465.47 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M736.7 55.72 L713.58 85.72 L734.9 109.46 L766.15 92.92 L766.51 84.35 L736.7 55.72 Z"
      /><path d="M736.7 55.72 L713.58 85.72 L734.9 109.46 L766.15 92.92 L766.51 84.35 L736.7 55.72 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1825.4 934.44 L1839.33 961.89 L1826.09 986.92 L1792.27 992.16 L1783.37 949.91 L1806.26 928.94 L1825.4 934.44 Z"
      /><path d="M1825.4 934.44 L1839.33 961.89 L1826.09 986.92 L1792.27 992.16 L1783.37 949.91 L1806.26 928.94 L1825.4 934.44 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M169.6 703.49 L168.41 703.39 L144.66 735.18 L156.91 761.78 L159.68 762.89 L192.91 741.55 L169.6 703.49 Z"
      /><path d="M169.6 703.49 L168.41 703.39 L144.66 735.18 L156.91 761.78 L159.68 762.89 L192.91 741.55 L169.6 703.49 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1494.58 416.59 L1459.28 381.03 L1438.49 421.87 L1444.3101 437.91 L1453.72 440.9 L1493.74 425.22 L1494.96 423.23 L1494.58 416.59 Z"
      /><path d="M1494.58 416.59 L1459.28 381.03 L1438.49 421.87 L1444.3101 437.91 L1453.72 440.9 L1493.74 425.22 L1494.96 423.23 L1494.58 416.59 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M453.65 266.38 L480.97 274.71 L484.25 299.79 L469.37 317.29 L468.69 317.27 L433.6 284.63 L453.65 266.38 Z"
      /><path d="M453.65 266.38 L480.97 274.71 L484.25 299.79 L469.37 317.29 L468.69 317.27 L433.6 284.63 L453.65 266.38 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1424.1 1028.36 L1392.4399 1050.62 L1373.8 1035.29 L1381 995.82 L1400.78 984.7 L1424.1 1028.36 Z"
      /><path d="M1424.1 1028.36 L1392.4399 1050.62 L1373.8 1035.29 L1381 995.82 L1400.78 984.7 L1424.1 1028.36 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M70.28 215.32 L51.94 252.8 L28.48 236.53 L30.86 206.87 L38.77 201.36 L70.28 215.32 Z"
      /><path d="M70.28 215.32 L51.94 252.8 L28.48 236.53 L30.86 206.87 L38.77 201.36 L70.28 215.32 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M761.96 637.96 L759.06 637.67 L740.09 652.32 L739.87 699.1 L757.95 703.32 L783.58 687.58 L787.13 665.4 L761.96 637.96 Z"
      /><path d="M761.96 637.96 L759.06 637.67 L740.09 652.32 L739.87 699.1 L757.95 703.32 L783.58 687.58 L787.13 665.4 L761.96 637.96 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M591.61 424.59 L606.03 443.03 L576.22 474.94 L574.44 474.38 L553.65 436.87 L553.73 436.71 L591.61 424.59 Z"
      /><path d="M591.61 424.59 L606.03 443.03 L576.22 474.94 L574.44 474.38 L553.65 436.87 L553.73 436.71 L591.61 424.59 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1682.8101 257.5 L1644.85 246.27 L1624.54 259.1 L1625.61 287.58 L1659.65 306.49 L1686.13 263.57 L1682.8101 257.5 Z"
      /><path d="M1682.8101 257.5 L1644.85 246.27 L1624.54 259.1 L1625.61 287.58 L1659.65 306.49 L1686.13 263.57 L1682.8101 257.5 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1343.6899 900.13 L1372.73 903.18 L1385.63 920.86 L1377.4399 943.06 L1342.6801 953.44 L1333.96 948.61 L1326.5601 922.09 L1343.6899 900.13 Z"
      /><path d="M1343.6899 900.13 L1372.73 903.18 L1385.63 920.86 L1377.4399 943.06 L1342.6801 953.44 L1333.96 948.61 L1326.5601 922.09 L1343.6899 900.13 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M367.9 0 L360.15 35.1 L316.26 44.51 L315.16 43.76 L309.2 0 L367.9 0 Z"
      /><path d="M367.9 0 L360.15 35.1 L316.26 44.51 L315.16 43.76 L309.2 0 L367.9 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1107.65 595.4 L1102.33 619.32 L1099.2 621.85 L1063.46 621.71 L1044.1 592.7 L1048.9301 574.04 L1066.76 568.26 L1107.65 595.4 Z"
      /><path d="M1107.65 595.4 L1102.33 619.32 L1099.2 621.85 L1063.46 621.71 L1044.1 592.7 L1048.9301 574.04 L1066.76 568.26 L1107.65 595.4 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1166.71 383.8 L1147.9301 382.35 L1117.8199 411.87 L1126.67 433.27 L1160.48 442.07 L1185.5699 413.55 L1166.71 383.8 Z"
      /><path d="M1166.71 383.8 L1147.9301 382.35 L1117.8199 411.87 L1126.67 433.27 L1160.48 442.07 L1185.5699 413.55 L1166.71 383.8 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1705.15 270.66 L1686.13 263.57 L1659.65 306.49 L1659.8101 307.07 L1703.45 330.84 L1723.52 308.33 L1705.15 270.66 Z"
      /><path d="M1705.15 270.66 L1686.13 263.57 L1659.65 306.49 L1659.8101 307.07 L1703.45 330.84 L1723.52 308.33 L1705.15 270.66 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1806.29 344.29 L1790.3101 331.65 L1766.95 335.08 L1742.8 376.59 L1742.84 378.24 L1747.1 385.24 L1800.54 395.43 L1803.25 393.57 L1806.29 344.29 Z"
      /><path d="M1806.29 344.29 L1790.3101 331.65 L1766.95 335.08 L1742.8 376.59 L1742.84 378.24 L1747.1 385.24 L1800.54 395.43 L1803.25 393.57 L1806.29 344.29 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1285.98 551.75 L1320.98 582.33 L1320.11 591.87 L1296.55 606.25 L1277.4301 594.26 L1276.86 561.7 L1285.98 551.75 Z"
      /><path d="M1285.98 551.75 L1320.98 582.33 L1320.11 591.87 L1296.55 606.25 L1277.4301 594.26 L1276.86 561.7 L1285.98 551.75 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M833.67 142.6 L815.31 122.68 L783.82 144.85 L790.08 158.31 L829.16 165.32 L833.67 142.6 Z"
      /><path d="M833.67 142.6 L815.31 122.68 L783.82 144.85 L790.08 158.31 L829.16 165.32 L833.67 142.6 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1333.96 948.61 L1303.7 964.98 L1311.08 1001.67 L1333.67 1003.58 L1349.42 988.6 L1342.6801 953.44 L1333.96 948.61 Z"
      /><path d="M1333.96 948.61 L1303.7 964.98 L1311.08 1001.67 L1333.67 1003.58 L1349.42 988.6 L1342.6801 953.44 L1333.96 948.61 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M325.44 965.51 L295.06 983.73 L288.96 1022.34 L358.19 1034.9 L359.46 1033.09 L357.18 990.02 L325.44 965.51 Z"
      /><path d="M325.44 965.51 L295.06 983.73 L288.96 1022.34 L358.19 1034.9 L359.46 1033.09 L357.18 990.02 L325.44 965.51 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M628.91 476.75 L632.75 480.01 L632.24 506.24 L605.5 519.91 L588.26 504.44 L587.43 489.04 L628.91 476.75 Z"
      /><path d="M628.91 476.75 L632.75 480.01 L632.24 506.24 L605.5 519.91 L588.26 504.44 L587.43 489.04 L628.91 476.75 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1457.87 871.73 L1478.34 909.48 L1462.87 928.99 L1437.28 933.22 L1418.38 916.55 L1426.4399 872.21 L1431.71 868.3 L1457.87 871.73 Z"
      /><path d="M1457.87 871.73 L1478.34 909.48 L1462.87 928.99 L1437.28 933.22 L1418.38 916.55 L1426.4399 872.21 L1431.71 868.3 L1457.87 871.73 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1920 700.6 L1871.98 704 L1872.36 751.89 L1920 759.3 L1920 700.6 Z"
      /><path d="M1920 700.6 L1871.98 704 L1872.36 751.89 L1920 759.3 L1920 700.6 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M221.03 494.45 L205.17 530.29 L207.19 534.83 L237.78 535.28 L244.34 502.07 L221.03 494.45 Z"
      /><path d="M221.03 494.45 L205.17 530.29 L207.19 534.83 L237.78 535.28 L244.34 502.07 L221.03 494.45 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M989.9 329.61 L972.22 297.47 L944.58 302.65 L934.04 334.2 L972.85 354.65 L989.9 329.61 Z"
      /><path d="M989.9 329.61 L972.22 297.47 L944.58 302.65 L934.04 334.2 L972.85 354.65 L989.9 329.61 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1366.34 725.41 L1342.1 736.29 L1356 772.05 L1391.6 774.3 L1398.35 750.09 L1366.34 725.41 Z"
      /><path d="M1366.34 725.41 L1342.1 736.29 L1356 772.05 L1391.6 774.3 L1398.35 750.09 L1366.34 725.41 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1239.04 704.5 L1255.1801 726.95 L1250.1801 735.56 L1216.34 748 L1198.74 729.21 L1214.1 706.66 L1239.04 704.5 Z"
      /><path d="M1239.04 704.5 L1255.1801 726.95 L1250.1801 735.56 L1216.34 748 L1198.74 729.21 L1214.1 706.66 L1239.04 704.5 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M975.02 89.76 L1010.44 94.13 L1022.56 109.96 L1017.44 136.34 L1001.79 146.38 L959.39 135.15 L975.02 89.76 Z"
      /><path d="M975.02 89.76 L1010.44 94.13 L1022.56 109.96 L1017.44 136.34 L1001.79 146.38 L959.39 135.15 L975.02 89.76 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M913.56 420.96 L938.12 440.17 L936.24 471.47 L912.11 485.86 L872.73 446.1 L874.91 434.17 L913.56 420.96 Z"
      /><path d="M913.56 420.96 L938.12 440.17 L936.24 471.47 L912.11 485.86 L872.73 446.1 L874.91 434.17 L913.56 420.96 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M644.71 890.79 L636.49 883.97 L603.56 889.34 L597.36 898.92 L611.45 939.11 L634.69 937.7 L649.86 919.29 L644.71 890.79 Z"
      /><path d="M644.71 890.79 L636.49 883.97 L603.56 889.34 L597.36 898.92 L611.45 939.11 L634.69 937.7 L649.86 919.29 L644.71 890.79 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1108.73 120.16 L1128.9399 134.34 L1129.22 162.93 L1089.84 179.95 L1064.64 160.66 L1079.65 126.4 L1108.73 120.16 Z"
      /><path d="M1108.73 120.16 L1128.9399 134.34 L1129.22 162.93 L1089.84 179.95 L1064.64 160.66 L1079.65 126.4 L1108.73 120.16 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M480.4 131.57 L487.93 174.64 L482.01 181.42 L456.13 184.28 L438.35 161.08 L459.41 125.18 L480.4 131.57 Z"
      /><path d="M480.4 131.57 L487.93 174.64 L482.01 181.42 L456.13 184.28 L438.35 161.08 L459.41 125.18 L480.4 131.57 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M695.36 575.01 L683.86 608.36 L669.14 610 L654.51 577.36 L671.28 558.67 L695.36 575.01 Z"
      /><path d="M695.36 575.01 L683.86 608.36 L669.14 610 L654.51 577.36 L671.28 558.67 L695.36 575.01 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M673.8 376.15 L627.61 378.97 L624.16 388.12 L645.17 426.9 L657.75 428.66 L677.49 415.18 L681.7 388.01 L673.8 376.15 Z"
      /><path d="M673.8 376.15 L627.61 378.97 L624.16 388.12 L645.17 426.9 L657.75 428.66 L677.49 415.18 L681.7 388.01 L673.8 376.15 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1250.1801 735.56 L1258.17 771.4 L1243.64 783.21 L1216.03 763.56 L1216.34 748 L1250.1801 735.56 Z"
      /><path d="M1250.1801 735.56 L1258.17 771.4 L1243.64 783.21 L1216.03 763.56 L1216.34 748 L1250.1801 735.56 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M424.82 336.66 L406.71 337.52 L387.03 356.63 L395.18 387.43 L422.51 386.7 L439.12 360.82 L431.35 340.3 L424.82 336.66 Z"
      /><path d="M424.82 336.66 L406.71 337.52 L387.03 356.63 L395.18 387.43 L422.51 386.7 L439.12 360.82 L431.35 340.3 L424.82 336.66 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M55.14 947.88 L44 926.65 L0 927 L0 975.8 L46.17 974.8 L55.14 947.88 Z"
      /><path d="M55.14 947.88 L44 926.65 L0 927 L0 975.8 L46.17 974.8 L55.14 947.88 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1331.91 531.87 L1342.1801 559.61 L1320.98 582.33 L1285.98 551.75 L1286.72 547.47 L1331.91 531.87 Z"
      /><path d="M1331.91 531.87 L1342.1801 559.61 L1320.98 582.33 L1285.98 551.75 L1286.72 547.47 L1331.91 531.87 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M659.57 209.16 L634.3 237.31 L614.82 221.7 L616.83 198.8 L649.11 195.35 L659.57 209.16 Z"
      /><path d="M659.57 209.16 L634.3 237.31 L614.82 221.7 L616.83 198.8 L649.11 195.35 L659.57 209.16 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M576.22 474.94 L574.44 474.38 L541 489.5 L541.1 512.38 L560.5 523.59 L588.26 504.44 L587.43 489.04 L576.22 474.94 Z"
      /><path d="M576.22 474.94 L574.44 474.38 L541 489.5 L541.1 512.38 L560.5 523.59 L588.26 504.44 L587.43 489.04 L576.22 474.94 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M183.88 559.66 L164.51 551.15 L143.49 572.87 L168.17 600.87 L180.01 594.82 L183.88 559.66 Z"
      /><path d="M183.88 559.66 L164.51 551.15 L143.49 572.87 L168.17 600.87 L180.01 594.82 L183.88 559.66 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M625.07 549.59 L605.73 532.69 L578.67 553.44 L583.21 565.78 L622.9 572.93 L625.07 549.59 Z"
      /><path d="M625.07 549.59 L605.73 532.69 L578.67 553.44 L583.21 565.78 L622.9 572.93 L625.07 549.59 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1089.5 528.79 L1044.89 502.75 L1042.7 503.74 L1023.8 549.93 L1048.9301 574.04 L1066.76 568.26 L1089.5 528.79 Z"
      /><path d="M1089.5 528.79 L1044.89 502.75 L1042.7 503.74 L1023.8 549.93 L1048.9301 574.04 L1066.76 568.26 L1089.5 528.79 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1260.28 1022.35 L1295.29 1039.72 L1278.6899 1071.14 L1243.16 1038.62 L1260.28 1022.35 Z"
      /><path d="M1260.28 1022.35 L1295.29 1039.72 L1278.6899 1071.14 L1243.16 1038.62 L1260.28 1022.35 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M104.42 636.37 L124.78 637.59 L133.73 655.33 L111.16 679.68 L85.62 663.37 L104.42 636.37 Z"
      /><path d="M104.42 636.37 L124.78 637.59 L133.73 655.33 L111.16 679.68 L85.62 663.37 L104.42 636.37 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M825.18 781.71 L838.73 793.09 L841.43 814.2 L821.69 842.89 L807.17 841.91 L784.79 801.16 L789.63 788.62 L825.18 781.71 Z"
      /><path d="M825.18 781.71 L838.73 793.09 L841.43 814.2 L821.69 842.89 L807.17 841.91 L784.79 801.16 L789.63 788.62 L825.18 781.71 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1486.66 601.61 L1477.99 642.06 L1433.1 642.15 L1423.52 626.58 L1447.5601 592.15 L1466.65 588.2 L1486.66 601.61 Z"
      /><path d="M1486.66 601.61 L1477.99 642.06 L1433.1 642.15 L1423.52 626.58 L1447.5601 592.15 L1466.65 588.2 L1486.66 601.61 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1748.7 144.97 L1791.05 181.08 L1734.89 208.17 L1721.6 164.96 L1748.7 144.97 Z"
      /><path d="M1748.7 144.97 L1791.05 181.08 L1734.89 208.17 L1721.6 164.96 L1748.7 144.97 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M764.33 575.07 L737.16 599.01 L759.06 637.67 L761.96 637.96 L795.29 610.68 L791.61 578.53 L764.33 575.07 Z"
      /><path d="M764.33 575.07 L737.16 599.01 L759.06 637.67 L761.96 637.96 L795.29 610.68 L791.61 578.53 L764.33 575.07 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M156.76 525.29 L164.51 551.15 L143.49 572.87 L129.31 572.72 L123.87 565.17 L125.66 538.84 L154.7 525.13 L156.76 525.29 Z"
      /><path d="M156.76 525.29 L164.51 551.15 L143.49 572.87 L129.31 572.72 L123.87 565.17 L125.66 538.84 L154.7 525.13 L156.76 525.29 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1632.8199 605.32 L1590.83 626.53 L1587.48 645.32 L1621.87 663.8 L1647.38 652.72 L1639.47 607.83 L1632.8199 605.32 Z"
      /><path d="M1632.8199 605.32 L1590.83 626.53 L1587.48 645.32 L1621.87 663.8 L1647.38 652.72 L1639.47 607.83 L1632.8199 605.32 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M310.76 729.02 L286.21 757.11 L323.42 784.99 L350.73 759.7 L351.05 747.2 L310.76 729.02 Z"
      /><path d="M310.76 729.02 L286.21 757.11 L323.42 784.99 L350.73 759.7 L351.05 747.2 L310.76 729.02 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M610.54 669.6 L651.03 673 L656.87 700.93 L610.68 703.98 L610.52 669.61 L610.54 669.6 Z"
      /><path d="M610.54 669.6 L651.03 673 L656.87 700.93 L610.68 703.98 L610.52 669.61 L610.54 669.6 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M153.48 60.47 L171.93 65.17 L187.92 111.21 L181.95 120.71 L150.18 128.19 L137.25 120.36 L133.46 81.79 L153.48 60.47 Z"
      /><path d="M153.48 60.47 L171.93 65.17 L187.92 111.21 L181.95 120.71 L150.18 128.19 L137.25 120.36 L133.46 81.79 L153.48 60.47 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M894.81 254.37 L917.6 274.59 L885.38 311.33 L862.79 302.24 L856.18 266.75 L894.81 254.37 Z"
      /><path d="M894.81 254.37 L917.6 274.59 L885.38 311.33 L862.79 302.24 L856.18 266.75 L894.81 254.37 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1178.4301 990.89 L1165.23 987.42 L1135.29 1002.51 L1147.22 1037.3199 L1168.14 1038.9301 L1179.35 992.63 L1178.4301 990.89 Z"
      /><path d="M1178.4301 990.89 L1165.23 987.42 L1135.29 1002.51 L1147.22 1037.3199 L1168.14 1038.9301 L1179.35 992.63 L1178.4301 990.89 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1437.89 795.58 L1391.86 774.86 L1380.27 823.74 L1426 826.41 L1438.87 810.08 L1437.89 795.58 Z"
      /><path d="M1437.89 795.58 L1391.86 774.86 L1380.27 823.74 L1426 826.41 L1438.87 810.08 L1437.89 795.58 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M732.54 412.78 L720 385.76 L681.7 388.01 L677.49 415.18 L709.1 432.51 L732.54 412.78 Z"
      /><path d="M732.54 412.78 L720 385.76 L681.7 388.01 L677.49 415.18 L709.1 432.51 L732.54 412.78 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M89.08 368.52 L94.43 369.47 L123.88 412.87 L116.79 424.3 L85.3 433.9 L74.18 426.98 L68.52 391.71 L89.08 368.52 Z"
      /><path d="M89.08 368.52 L94.43 369.47 L123.88 412.87 L116.79 424.3 L85.3 433.9 L74.18 426.98 L68.52 391.71 L89.08 368.52 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1533.77 641.08 L1489.5601 657.08 L1489.09 667.11 L1516.39 697.18 L1540.0699 684.66 L1542.27 649.24 L1533.77 641.08 Z"
      /><path d="M1533.77 641.08 L1489.5601 657.08 L1489.09 667.11 L1516.39 697.18 L1540.0699 684.66 L1542.27 649.24 L1533.77 641.08 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1173.0699 35.97 L1137.3199 62.67 L1165.5699 97.6 L1200.3101 83.52 L1200.78 52.4 L1173.0699 35.97 Z"
      /><path d="M1173.0699 35.97 L1137.3199 62.67 L1165.5699 97.6 L1200.3101 83.52 L1200.78 52.4 L1173.0699 35.97 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1307.26 269.82 L1315.33 271.52 L1324.33 307.61 L1308.17 327.93 L1274.03 318.52 L1269.62 298.37 L1307.26 269.82 Z"
      /><path d="M1307.26 269.82 L1315.33 271.52 L1324.33 307.61 L1308.17 327.93 L1274.03 318.52 L1269.62 298.37 L1307.26 269.82 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1259.03 66.54 L1222.41 100.04 L1226.0699 115.48 L1249.65 129.63 L1285.26 93.47 L1283.64 85.19 L1259.03 66.54 Z"
      /><path d="M1259.03 66.54 L1222.41 100.04 L1226.0699 115.48 L1249.65 129.63 L1285.26 93.47 L1283.64 85.19 L1259.03 66.54 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1081.6801 989.5 L1114.84 990.79 L1120.85 998.52 L1102.59 1034.1899 L1082.08 1036.97 L1074.35 1030.89 L1081.6801 989.5 Z"
      /><path d="M1081.6801 989.5 L1114.84 990.79 L1120.85 998.52 L1102.59 1034.1899 L1082.08 1036.97 L1074.35 1030.89 L1081.6801 989.5 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1920 894.5 L1920 841.1 L1883.42 848.34 L1877.5699 887.77 L1920 894.5 Z"
      /><path d="M1920 894.5 L1920 841.1 L1883.42 848.34 L1877.5699 887.77 L1920 894.5 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M937.97 792.54 L976.93 816.13 L968.72 838.72 L932.61 839.71 L922.21 809.48 L937.97 792.54 Z"
      /><path d="M937.97 792.54 L976.93 816.13 L968.72 838.72 L932.61 839.71 L922.21 809.48 L937.97 792.54 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M125.76 773.69 L119.69 804.35 L99.61 809.61 L85.23 799.7 L87.57 760.52 L105.54 755.78 L125.76 773.69 Z"
      /><path d="M125.76 773.69 L119.69 804.35 L99.61 809.61 L85.23 799.7 L87.57 760.52 L105.54 755.78 L125.76 773.69 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1272.59 517.93 L1254.5 484.83 L1223.7 488.04 L1213.23 513.76 L1233.73 533.47 L1272.52 518.23 L1272.59 517.93 Z"
      /><path d="M1272.59 517.93 L1254.5 484.83 L1223.7 488.04 L1213.23 513.76 L1233.73 533.47 L1272.52 518.23 L1272.59 517.93 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1656.27 706.76 L1630.04 717.57 L1627.83 727.63 L1648.48 763.49 L1695.37 741.63 L1696.33 732.66 L1656.27 706.76 Z"
      /><path d="M1656.27 706.76 L1630.04 717.57 L1627.83 727.63 L1648.48 763.49 L1695.37 741.63 L1696.33 732.66 L1656.27 706.76 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1189.92 291.1 L1175.36 334.49 L1140.51 328.02 L1155.96 288.74 L1189.92 291.1 Z"
      /><path d="M1189.92 291.1 L1175.36 334.49 L1140.51 328.02 L1155.96 288.74 L1189.92 291.1 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M126.47 231.31 L111.83 234.5 L92.84 267.22 L104.94 298.43 L121.68 302.89 L155.2 281.85 L151.41 246.97 L126.47 231.31 Z"
      /><path d="M126.47 231.31 L111.83 234.5 L92.84 267.22 L104.94 298.43 L121.68 302.89 L155.2 281.85 L151.41 246.97 L126.47 231.31 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M957 136.4 L930.18 131.54 L901.98 163.58 L928.41 202.01 L932.66 202.83 L955.41 186.63 L957 136.4 Z"
      /><path d="M957 136.4 L930.18 131.54 L901.98 163.58 L928.41 202.01 L932.66 202.83 L955.41 186.63 L957 136.4 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M225.26 339.52 L236.45 382.13 L215.59 404.28 L192.2 387.02 L196.63 340.12 L221.27 336.96 L225.26 339.52 Z"
      /><path d="M225.26 339.52 L236.45 382.13 L215.59 404.28 L192.2 387.02 L196.63 340.12 L221.27 336.96 L225.26 339.52 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M583.21 565.78 L622.9 572.93 L626.12 578.99 L625.73 580.36 L599.07 602.77 L575.39 590.19 L583.21 565.78 Z"
      /><path d="M583.21 565.78 L622.9 572.93 L626.12 578.99 L625.73 580.36 L599.07 602.77 L575.39 590.19 L583.21 565.78 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M775.58 103.82 L814.17 105.57 L815.31 122.68 L783.82 144.85 L772.63 139.14 L775.58 103.82 Z"
      /><path d="M775.58 103.82 L814.17 105.57 L815.31 122.68 L783.82 144.85 L772.63 139.14 L775.58 103.82 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1839.33 961.89 L1871.77 962.79 L1883.04 988.7 L1857.67 1020.59 L1852.9 1020.41 L1826.09 986.92 L1839.33 961.89 Z"
      /><path d="M1839.33 961.89 L1871.77 962.79 L1883.04 988.7 L1857.67 1020.59 L1852.9 1020.41 L1826.09 986.92 L1839.33 961.89 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1355 0 L1355 2.45 L1373.36 37.18 L1397.16 43.26 L1432.09 0.23 L1432.1 0 L1355 0 Z"
      /><path d="M1355 0 L1355 2.45 L1373.36 37.18 L1397.16 43.26 L1432.09 0.23 L1432.1 0 L1355 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1277.67 948.72 L1249.76 941.95 L1228.23 965.84 L1237.03 985.87 L1261.96 994.31 L1282.98 958.18 L1277.67 948.72 Z"
      /><path d="M1277.67 948.72 L1249.76 941.95 L1228.23 965.84 L1237.03 985.87 L1261.96 994.31 L1282.98 958.18 L1277.67 948.72 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1297.21 1038.64 L1334.95 1052.67 L1336.5 1080 L1278.8 1080 L1278.6899 1071.14 L1295.29 1039.72 L1297.21 1038.64 Z"
      /><path d="M1297.21 1038.64 L1334.95 1052.67 L1336.5 1080 L1278.8 1080 L1278.6899 1071.14 L1295.29 1039.72 L1297.21 1038.64 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M322.6 534.97 L301.9 507.45 L276.79 517.99 L271.98 541.35 L289.71 557.58 L322.6 534.97 Z"
      /><path d="M322.6 534.97 L301.9 507.45 L276.79 517.99 L271.98 541.35 L289.71 557.58 L322.6 534.97 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M313.5 448.11 L280.83 439.21 L263.72 465.47 L265.48 471.98 L306.12 488.08 L317.71 478.3 L313.5 448.11 Z"
      /><path d="M313.5 448.11 L280.83 439.21 L263.72 465.47 L265.48 471.98 L306.12 488.08 L317.71 478.3 L313.5 448.11 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1875.01 228.34 L1870.62 287.28 L1848.23 292.33 L1825.05 279.94 L1821.25 232.97 L1861.79 218.72 L1875.01 228.34 Z"
      /><path d="M1875.01 228.34 L1870.62 287.28 L1848.23 292.33 L1825.05 279.94 L1821.25 232.97 L1861.79 218.72 L1875.01 228.34 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M39.72 514.88 L51.32 547.29 L38.41 559.12 L0.92 537.07 L35.48 513.66 L39.72 514.88 Z"
      /><path d="M39.72 514.88 L51.32 547.29 L38.41 559.12 L0.92 537.07 L35.48 513.66 L39.72 514.88 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M838.52 884.17 L879.04 890.19 L879.52 890.79 L881.11 913.5 L857.45 938.57 L842.5 934.86 L826.23 901.28 L838.52 884.17 Z"
      /><path d="M838.52 884.17 L879.04 890.19 L879.52 890.79 L881.11 913.5 L857.45 938.57 L842.5 934.86 L826.23 901.28 L838.52 884.17 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1060.09 869.56 L1041.4 893.66 L1041.86 895.96 L1067.77 922.53 L1084.63 923.49 L1096.52 907.91 L1086.1 874.92 L1060.09 869.56 Z"
      /><path d="M1060.09 869.56 L1041.4 893.66 L1041.86 895.96 L1067.77 922.53 L1084.63 923.49 L1096.52 907.91 L1086.1 874.92 L1060.09 869.56 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1316.11 206.44 L1299.5 175.74 L1259.36 186.73 L1257.5699 201.83 L1284.3101 227.04 L1316.11 206.44 Z"
      /><path d="M1316.11 206.44 L1299.5 175.74 L1259.36 186.73 L1257.5699 201.83 L1284.3101 227.04 L1316.11 206.44 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M670.24 1004.04 L635.2 989.26 L633.99 989.74 L628.58 1029.45 L643.02 1035.6899 L670.31 1013.63 L670.24 1004.04 Z"
      /><path d="M670.24 1004.04 L635.2 989.26 L633.99 989.74 L628.58 1029.45 L643.02 1035.6899 L670.31 1013.63 L670.24 1004.04 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M928.41 202.01 L932.66 202.83 L952.17 241.84 L917.95 274.61 L917.6 274.59 L894.81 254.37 L894.37 223.33 L928.41 202.01 Z"
      /><path d="M928.41 202.01 L932.66 202.83 L952.17 241.84 L917.95 274.61 L917.6 274.59 L894.81 254.37 L894.37 223.33 L928.41 202.01 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1875.21 637.64 L1860.4301 694.84 L1841.14 696.19 L1804.1 649.95 L1809.28 636.85 L1870.65 633.44 L1875.21 637.64 Z"
      /><path d="M1875.21 637.64 L1860.4301 694.84 L1841.14 696.19 L1804.1 649.95 L1809.28 636.85 L1870.65 633.44 L1875.21 637.64 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1001.39 996.75 L966.98 991.76 L958.73 1028.3101 L983.58 1045.48 L1002.39 1031.47 L1001.39 996.75 Z"
      /><path d="M1001.39 996.75 L966.98 991.76 L958.73 1028.3101 L983.58 1045.48 L1002.39 1031.47 L1001.39 996.75 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M532.67 447.06 L503.77 428.49 L486.48 437.54 L482.72 447.92 L509.55 477.17 L523.72 474.55 L532.67 447.06 Z"
      /><path d="M532.67 447.06 L503.77 428.49 L486.48 437.54 L482.72 447.92 L509.55 477.17 L523.72 474.55 L532.67 447.06 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M200.98 553.18 L216.25 569.85 L204.59 599.81 L180.01 594.82 L183.88 559.66 L200.98 553.18 Z"
      /><path d="M200.98 553.18 L216.25 569.85 L204.59 599.81 L180.01 594.82 L183.88 559.66 L200.98 553.18 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1286.72 547.47 L1272.52 518.23 L1233.73 533.47 L1231.6801 561.6 L1237.75 565.78 L1276.86 561.7 L1285.98 551.75 L1286.72 547.47 Z"
      /><path d="M1286.72 547.47 L1272.52 518.23 L1233.73 533.47 L1231.6801 561.6 L1237.75 565.78 L1276.86 561.7 L1285.98 551.75 L1286.72 547.47 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1837.28 337.23 L1806.29 344.29 L1803.25 393.57 L1835.27 398.19 L1864.6 370.36 L1865.73 359.89 L1837.28 337.23 Z"
      /><path d="M1837.28 337.23 L1806.29 344.29 L1803.25 393.57 L1835.27 398.19 L1864.6 370.36 L1865.73 359.89 L1837.28 337.23 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M358.13 347.46 L387.03 356.63 L395.18 387.43 L386.27 398.57 L346.18 392.15 L340.74 376.24 L354.79 348.54 L358.13 347.46 Z"
      /><path d="M358.13 347.46 L387.03 356.63 L395.18 387.43 L386.27 398.57 L346.18 392.15 L340.74 376.24 L354.79 348.54 L358.13 347.46 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1200.14 201.37 L1230.11 220.28 L1230.21 248.09 L1196.38 259.35 L1176.76 241.35 L1175.3199 222.58 L1200.14 201.37 Z"
      /><path d="M1200.14 201.37 L1230.11 220.28 L1230.21 248.09 L1196.38 259.35 L1176.76 241.35 L1175.3199 222.58 L1200.14 201.37 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M610.52 669.61 L585.45 662.54 L556.45 692.3 L556.73 695.47 L602.21 715.47 L610.68 703.98 L610.52 669.61 Z"
      /><path d="M610.52 669.61 L585.45 662.54 L556.45 692.3 L556.73 695.47 L602.21 715.47 L610.68 703.98 L610.52 669.61 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M204.34 47.76 L221.2 55.86 L228.9 100.96 L187.92 111.21 L171.93 65.17 L204.34 47.76 Z"
      /><path d="M204.34 47.76 L221.2 55.86 L228.9 100.96 L187.92 111.21 L171.93 65.17 L204.34 47.76 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M276.79 517.99 L271.98 541.35 L248.3 546.83 L237.78 535.28 L244.34 502.07 L253.38 498.8 L276.79 517.99 Z"
      /><path d="M276.79 517.99 L271.98 541.35 L248.3 546.83 L237.78 535.28 L244.34 502.07 L253.38 498.8 L276.79 517.99 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1392.4399 1050.62 L1393.7 1080 L1336.5 1080 L1334.95 1052.67 L1346.4301 1038.15 L1373.8 1035.29 L1392.4399 1050.62 Z"
      /><path d="M1392.4399 1050.62 L1393.7 1080 L1336.5 1080 L1334.95 1052.67 L1346.4301 1038.15 L1373.8 1035.29 L1392.4399 1050.62 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1386.0699 868.1 L1372.73 903.18 L1343.6899 900.13 L1329.34 865.52 L1375.4399 852.93 L1386.0699 868.1 Z"
      /><path d="M1386.0699 868.1 L1372.73 903.18 L1343.6899 900.13 L1329.34 865.52 L1375.4399 852.93 L1386.0699 868.1 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1649.03 433.26 L1620.51 405.76 L1596.2 432.19 L1596.64 433.25 L1629.22 450.47 L1649.01 439 L1649.03 433.26 Z"
      /><path d="M1649.03 433.26 L1620.51 405.76 L1596.2 432.19 L1596.64 433.25 L1629.22 450.47 L1649.01 439 L1649.03 433.26 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M655.9 294.31 L698.14 295.6 L700.69 307.47 L677.02 341.68 L656.1 330.73 L655.9 294.31 Z"
      /><path d="M655.9 294.31 L698.14 295.6 L700.69 307.47 L677.02 341.68 L656.1 330.73 L655.9 294.31 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M368.32 727.8 L382.83 728.75 L413.76 752.58 L417.28 767.92 L386.01 792.03 L350.73 759.7 L351.05 747.2 L368.32 727.8 Z"
      /><path d="M368.32 727.8 L382.83 728.75 L413.76 752.58 L417.28 767.92 L386.01 792.03 L350.73 759.7 L351.05 747.2 L368.32 727.8 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1020.96 927.31 L1030.2 946.16 L1007.98 964.05 L988.39 954.11 L983.47 939.39 L1000.13 920.84 L1020.96 927.31 Z"
      /><path d="M1020.96 927.31 L1030.2 946.16 L1007.98 964.05 L988.39 954.11 L983.47 939.39 L1000.13 920.84 L1020.96 927.31 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M693.22 855.86 L684.07 842.62 L641.24 851.76 L636.49 883.97 L644.71 890.79 L684.8 881.69 L693.22 855.86 Z"
      /><path d="M693.22 855.86 L684.07 842.62 L641.24 851.76 L636.49 883.97 L644.71 890.79 L684.8 881.69 L693.22 855.86 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1283.85 894.29 L1268.97 868.47 L1227.04 871.53 L1226.24 907.47 L1239.89 915.02 L1283.78 895.05 L1283.85 894.29 Z"
      /><path d="M1283.85 894.29 L1268.97 868.47 L1227.04 871.53 L1226.24 907.47 L1239.89 915.02 L1283.78 895.05 L1283.85 894.29 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M824.03 628.74 L795.29 610.68 L761.96 637.96 L787.13 665.4 L818.62 653.73 L824.03 628.74 Z"
      /><path d="M824.03 628.74 L795.29 610.68 L761.96 637.96 L787.13 665.4 L818.62 653.73 L824.03 628.74 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1448.14 100.48 L1405.9399 98.43 L1406.36 137.63 L1418.35 145.5 L1457.83 117.45 L1448.14 100.48 Z"
      /><path d="M1448.14 100.48 L1405.9399 98.43 L1406.36 137.63 L1418.35 145.5 L1457.83 117.45 L1448.14 100.48 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M903.8 506.74 L845.17 497.66 L835.03 518.61 L849.66 546.38 L893.09 546.65 L908.74 529.58 L903.8 506.74 Z"
      /><path d="M903.8 506.74 L845.17 497.66 L835.03 518.61 L849.66 546.38 L893.09 546.65 L908.74 529.58 L903.8 506.74 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1128.03 344.74 L1147.9301 382.35 L1117.8199 411.87 L1103.05 405.39 L1091.98 373.07 L1111.92 347.33 L1128.03 344.74 Z"
      /><path d="M1128.03 344.74 L1147.9301 382.35 L1117.8199 411.87 L1103.05 405.39 L1091.98 373.07 L1111.92 347.33 L1128.03 344.74 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1313.46 782.43 L1326.7 732.88 L1289.79 743.38 L1284.02 773.12 L1297.38 787.42 L1313.46 782.43 Z"
      /><path d="M1313.46 782.43 L1326.7 732.88 L1289.79 743.38 L1284.02 773.12 L1297.38 787.42 L1313.46 782.43 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1277.4301 594.26 L1296.55 606.25 L1294.51 627.32 L1261.79 639.1 L1252.58 634.16 L1243.72 613.08 L1247.91 605.29 L1277.4301 594.26 Z"
      /><path d="M1277.4301 594.26 L1296.55 606.25 L1294.51 627.32 L1261.79 639.1 L1252.58 634.16 L1243.72 613.08 L1247.91 605.29 L1277.4301 594.26 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1079.65 126.4 L1064.64 160.66 L1056.55 162.49 L1017.44 136.34 L1022.56 109.96 L1058.45 102.17 L1079.65 126.4 Z"
      /><path d="M1079.65 126.4 L1064.64 160.66 L1056.55 162.49 L1017.44 136.34 L1022.56 109.96 L1058.45 102.17 L1079.65 126.4 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1294.51 627.32 L1313.95 648.22 L1310.23 661.36 L1278.47 676.99 L1272.05 674.12 L1261.79 639.1 L1294.51 627.32 Z"
      /><path d="M1294.51 627.32 L1313.95 648.22 L1310.23 661.36 L1278.47 676.99 L1272.05 674.12 L1261.79 639.1 L1294.51 627.32 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M28.48 236.53 L51.94 252.8 L54.22 261.12 L45.17 274.73 L0 272.9 L0 244.8 L28.48 236.53 Z"
      /><path d="M28.48 236.53 L51.94 252.8 L54.22 261.12 L45.17 274.73 L0 272.9 L0 244.8 L28.48 236.53 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1364.64 335.87 L1393.1 345.75 L1398.83 382.64 L1392.42 393.75 L1355.6801 389.41 L1346.84 357.43 L1364.64 335.87 Z"
      /><path d="M1364.64 335.87 L1393.1 345.75 L1398.83 382.64 L1392.42 393.75 L1355.6801 389.41 L1346.84 357.43 L1364.64 335.87 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M329.63 145.78 L347.28 154.79 L357.43 174.82 L348.85 200.54 L340.18 205.31 L314.55 193.93 L314.36 157.28 L328.7 145.89 L329.63 145.78 Z"
      /><path d="M329.63 145.78 L347.28 154.79 L357.43 174.82 L348.85 200.54 L340.18 205.31 L314.55 193.93 L314.36 157.28 L328.7 145.89 L329.63 145.78 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M982.78 734.49 L983.45 762.21 L939.1 779.31 L922.52 755.08 L944.61 727.04 L982.78 734.49 Z"
      /><path d="M982.78 734.49 L983.45 762.21 L939.1 779.31 L922.52 755.08 L944.61 727.04 L982.78 734.49 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M346.14 290.12 L320.97 323.75 L285.94 292.46 L298.77 263.69 L346.14 290.12 Z"
      /><path d="M346.14 290.12 L320.97 323.75 L285.94 292.46 L298.77 263.69 L346.14 290.12 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M674.46 211.8 L671.67 212.56 L669.94 254.08 L694.27 258.92 L699.26 253.72 L699.68 221.61 L674.46 211.8 Z"
      /><path d="M674.46 211.8 L671.67 212.56 L669.94 254.08 L694.27 258.92 L699.26 253.72 L699.68 221.61 L674.46 211.8 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M262.44 785.3 L254.85 786.24 L227.84 819.7 L240.95 841.26 L281.04 842.75 L287.2 816.13 L262.44 785.3 Z"
      /><path d="M262.44 785.3 L254.85 786.24 L227.84 819.7 L240.95 841.26 L281.04 842.75 L287.2 816.13 L262.44 785.3 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1226.24 907.47 L1212.9399 913.57 L1199.78 953.18 L1201.67 957.84 L1228.23 965.84 L1249.76 941.95 L1239.89 915.02 L1226.24 907.47 Z"
      /><path d="M1226.24 907.47 L1212.9399 913.57 L1199.78 953.18 L1201.67 957.84 L1228.23 965.84 L1249.76 941.95 L1239.89 915.02 L1226.24 907.47 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M0 202.7 L30.86 206.87 L28.48 236.53 L0 244.8 L0 202.7 Z"
      /><path d="M0 202.7 L30.86 206.87 L28.48 236.53 L0 244.8 L0 202.7 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M332.53 537.24 L322.6 534.97 L289.71 557.58 L290.11 574.14 L312.83 591.24 L342.17 573.17 L332.53 537.24 Z"
      /><path d="M332.53 537.24 L322.6 534.97 L289.71 557.58 L290.11 574.14 L312.83 591.24 L342.17 573.17 L332.53 537.24 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1696.63 450.35 L1720.85 493.59 L1717.42 497.01 L1687.22 506.56 L1658.9301 496.84 L1658.86 496.74 L1669.61 455.92 L1696.63 450.35 Z"
      /><path d="M1696.63 450.35 L1720.85 493.59 L1717.42 497.01 L1687.22 506.56 L1658.9301 496.84 L1658.86 496.74 L1669.61 455.92 L1696.63 450.35 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M328.7 145.89 L314.36 157.28 L278.91 151.42 L277.99 130.71 L301.14 106.97 L328.7 145.89 Z"
      /><path d="M328.7 145.89 L314.36 157.28 L278.91 151.42 L277.99 130.71 L301.14 106.97 L328.7 145.89 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M227.84 819.7 L240.95 841.26 L223.55 881.63 L220.47 883.01 L185.49 868.11 L180.3 855.2 L202.41 814.56 L227.84 819.7 Z"
      /><path d="M227.84 819.7 L240.95 841.26 L223.55 881.63 L220.47 883.01 L185.49 868.11 L180.3 855.2 L202.41 814.56 L227.84 819.7 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M621.76 640.02 L610.54 669.6 L651.03 673 L661.1 653.16 L658.71 648.64 L621.76 640.02 Z"
      /><path d="M621.76 640.02 L610.54 669.6 L651.03 673 L661.1 653.16 L658.71 648.64 L621.76 640.02 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M294.69 252.09 L248.71 245.48 L223.36 269.56 L223.3 270.05 L233.19 286.06 L272.56 299.59 L285.94 292.46 L298.77 263.69 L297.73 255.08 L294.69 252.09 Z"
      /><path d="M294.69 252.09 L248.71 245.48 L223.36 269.56 L223.3 270.05 L233.19 286.06 L272.56 299.59 L285.94 292.46 L298.77 263.69 L297.73 255.08 L294.69 252.09 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M289.71 557.58 L290.11 574.14 L262.99 589.74 L249.23 583.1 L241.26 569.85 L248.3 546.83 L271.98 541.35 L289.71 557.58 Z"
      /><path d="M289.71 557.58 L290.11 574.14 L262.99 589.74 L249.23 583.1 L241.26 569.85 L248.3 546.83 L271.98 541.35 L289.71 557.58 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M502.88 86.18 L504.47 119.59 L480.4 131.57 L459.41 125.18 L452.48 114.76 L469.53 70.69 L502.88 86.18 Z"
      /><path d="M502.88 86.18 L504.47 119.59 L480.4 131.57 L459.41 125.18 L452.48 114.76 L469.53 70.69 L502.88 86.18 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1099.2 621.85 L1063.46 621.71 L1043.42 652.95 L1044.83 662.1 L1089.38 673.18 L1093.29 670.76 L1099.2 621.85 Z"
      /><path d="M1099.2 621.85 L1063.46 621.71 L1043.42 652.95 L1044.83 662.1 L1089.38 673.18 L1093.29 670.76 L1099.2 621.85 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M204.59 599.81 L180.01 594.82 L168.17 600.87 L162.59 613 L177.38 644.64 L184.66 647.07 L219.42 626.68 L216.99 614.51 L204.59 599.81 Z"
      /><path d="M204.59 599.81 L180.01 594.82 L168.17 600.87 L162.59 613 L177.38 644.64 L184.66 647.07 L219.42 626.68 L216.99 614.51 L204.59 599.81 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M359.64 580.4 L342.17 573.17 L312.83 591.24 L312.53 608.53 L342.26 634.64 L352.01 635.46 L363.6 623.36 L359.64 580.4 Z"
      /><path d="M359.64 580.4 L342.17 573.17 L312.83 591.24 L312.53 608.53 L342.26 634.64 L352.01 635.46 L363.6 623.36 L359.64 580.4 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M536.15 192.35 L516.66 170.99 L487.93 174.64 L482.01 181.42 L498.24 224.93 L502.95 224.37 L535.58 198.25 L536.15 192.35 Z"
      /><path d="M536.15 192.35 L516.66 170.99 L487.93 174.64 L482.01 181.42 L498.24 224.93 L502.95 224.37 L535.58 198.25 L536.15 192.35 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M223.55 881.63 L269.44 896.61 L279.61 911.81 L253.69 952.19 L245.17 954.12 L211.35 923.47 L220.47 883.01 L223.55 881.63 Z"
      /><path d="M223.55 881.63 L269.44 896.61 L279.61 911.81 L253.69 952.19 L245.17 954.12 L211.35 923.47 L220.47 883.01 L223.55 881.63 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M664.9 0 L610.9 0 L609.89 33.14 L626.81 47.71 L665.33 33.02 L664.9 0 Z"
      /><path d="M664.9 0 L610.9 0 L609.89 33.14 L626.81 47.71 L665.33 33.02 L664.9 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1883.04 988.7 L1920 994.7 L1920 1032.5 L1877.12 1039.75 L1857.67 1020.59 L1883.04 988.7 Z"
      /><path d="M1883.04 988.7 L1920 994.7 L1920 1032.5 L1877.12 1039.75 L1857.67 1020.59 L1883.04 988.7 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M115.21 730.98 L105.54 755.78 L87.57 760.52 L69.73 751.45 L67.92 746.7 L81.73 712.01 L87.33 711.81 L115.21 730.98 Z"
      /><path d="M115.21 730.98 L105.54 755.78 L87.57 760.52 L69.73 751.45 L67.92 746.7 L81.73 712.01 L87.33 711.81 L115.21 730.98 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M374.04 110.31 L380.48 116.2 L376.64 135.05 L347.28 154.79 L329.63 145.78 L347.01 113.6 L374.04 110.31 Z"
      /><path d="M374.04 110.31 L380.48 116.2 L376.64 135.05 L347.28 154.79 L329.63 145.78 L347.01 113.6 L374.04 110.31 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1523.46 165.28 L1560.88 185.1 L1562.77 202.96 L1547.48 220.29 L1513.15 221 L1495.34 187.86 L1523.46 165.28 Z"
      /><path d="M1523.46 165.28 L1560.88 185.1 L1562.77 202.96 L1547.48 220.29 L1513.15 221 L1495.34 187.86 L1523.46 165.28 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1685.75 91.93 L1660.9301 101.88 L1649.3199 135.7 L1685.42 157.97 L1693.27 155.34 L1708.21 102.79 L1685.75 91.93 Z"
      /><path d="M1685.75 91.93 L1660.9301 101.88 L1649.3199 135.7 L1685.42 157.97 L1693.27 155.34 L1708.21 102.79 L1685.75 91.93 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M364.5 444.16 L332.83 426.99 L313.5 448.11 L317.71 478.3 L345.91 484.61 L366.76 467.25 L364.5 444.16 Z"
      /><path d="M364.5 444.16 L332.83 426.99 L313.5 448.11 L317.71 478.3 L345.91 484.61 L366.76 467.25 L364.5 444.16 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M664.09 707.68 L656.87 700.93 L610.68 703.98 L602.21 715.47 L604.66 738.71 L665.14 738.08 L664.09 707.68 Z"
      /><path d="M664.09 707.68 L656.87 700.93 L610.68 703.98 L602.21 715.47 L604.66 738.71 L665.14 738.08 L664.09 707.68 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1728.53 1004.45 L1731.23 1027.51 L1716.08 1045.41 L1682.91 1039.1801 L1674.46 1015.79 L1684.95 998.44 L1728.53 1004.45 Z"
      /><path d="M1728.53 1004.45 L1731.23 1027.51 L1716.08 1045.41 L1682.91 1039.1801 L1674.46 1015.79 L1684.95 998.44 L1728.53 1004.45 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1373.36 37.18 L1351.62 69.64 L1341.9 71.49 L1319 56.45 L1316.4 44.46 L1355 2.45 L1373.36 37.18 Z"
      /><path d="M1373.36 37.18 L1351.62 69.64 L1341.9 71.49 L1319 56.45 L1316.4 44.46 L1355 2.45 L1373.36 37.18 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1731.23 1027.51 L1770.08 1043.25 L1769.3 1080 L1720.1 1080 L1716.08 1045.41 L1731.23 1027.51 Z"
      /><path d="M1731.23 1027.51 L1770.08 1043.25 L1769.3 1080 L1720.1 1080 L1716.08 1045.41 L1731.23 1027.51 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M413.99 601.69 L442.38 605.9 L456.22 640.31 L451.38 650.76 L416.9 663.88 L398.99 621.76 L413.99 601.69 Z"
      /><path d="M413.99 601.69 L442.38 605.9 L456.22 640.31 L451.38 650.76 L416.9 663.88 L398.99 621.76 L413.99 601.69 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M418.06 1021.67 L438.25 1041.03 L438.3 1080 L358.6 1080 L358.19 1034.9 L359.46 1033.09 L418.06 1021.67 Z"
      /><path d="M418.06 1021.67 L438.25 1041.03 L438.3 1080 L358.6 1080 L358.19 1034.9 L359.46 1033.09 L418.06 1021.67 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M137.25 120.36 L150.18 128.19 L147.24 178.46 L138.53 182.88 L98.49 168.81 L97.36 132.02 L97.74 131.52 L137.25 120.36 Z"
      /><path d="M137.25 120.36 L150.18 128.19 L147.24 178.46 L138.53 182.88 L98.49 168.81 L97.36 132.02 L97.74 131.52 L137.25 120.36 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1351.62 69.64 L1341.9 71.49 L1331.58 107.63 L1346.24 123.13 L1362.1899 123.16 L1382.48 91.62 L1351.62 69.64 Z"
      /><path d="M1351.62 69.64 L1341.9 71.49 L1331.58 107.63 L1346.24 123.13 L1362.1899 123.16 L1382.48 91.62 L1351.62 69.64 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1748.97 660.26 L1729.78 626.92 L1704.73 628.04 L1677.38 663.45 L1721.23 700.74 L1748.97 660.26 Z"
      /><path d="M1748.97 660.26 L1729.78 626.92 L1704.73 628.04 L1677.38 663.45 L1721.23 700.74 L1748.97 660.26 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M55.45 991.36 L46.17 974.8 L0 975.8 L0 1020.1 L40.81 1025.8199 L55.45 991.36 Z"
      /><path d="M55.45 991.36 L46.17 974.8 L0 975.8 L0 1020.1 L40.81 1025.8199 L55.45 991.36 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M45.17 274.73 L0 272.9 L0 312.9 L35.12 316.65 L47.72 304.12 L45.17 274.73 Z"
      /><path d="M45.17 274.73 L0 272.9 L0 312.9 L35.12 316.65 L47.72 304.12 L45.17 274.73 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M396.22 168.86 L357.43 174.82 L348.85 200.54 L385.96 213.95 L402.33 197.04 L400.17 170.57 L396.22 168.86 Z"
      /><path d="M396.22 168.86 L357.43 174.82 L348.85 200.54 L385.96 213.95 L402.33 197.04 L400.17 170.57 L396.22 168.86 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M517.93 37.77 L527.47 47.56 L527.64 70.85 L502.88 86.18 L469.53 70.69 L466.45 64 L486.19 37.92 L517.93 37.77 Z"
      /><path d="M517.93 37.77 L527.47 47.56 L527.64 70.85 L502.88 86.18 L469.53 70.69 L466.45 64 L486.19 37.92 L517.93 37.77 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1767.3199 72.9 L1789.02 73.93 L1807.24 111.73 L1798.15 120.87 L1753.01 118.95 L1767.3199 72.9 Z"
      /><path d="M1767.3199 72.9 L1789.02 73.93 L1807.24 111.73 L1798.15 120.87 L1753.01 118.95 L1767.3199 72.9 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M128.51 698.36 L121.15 728.44 L115.21 730.98 L87.33 711.81 L112.05 684.53 L128.51 698.36 Z"
      /><path d="M128.51 698.36 L121.15 728.44 L115.21 730.98 L87.33 711.81 L112.05 684.53 L128.51 698.36 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1557.78 1024.0601 L1564.11 1029.52 L1558.5 1080 L1507 1080 L1505.8101 1037.59 L1522.37 1022.36 L1557.78 1024.0601 Z"
      /><path d="M1557.78 1024.0601 L1564.11 1029.52 L1558.5 1080 L1507 1080 L1505.8101 1037.59 L1522.37 1022.36 L1557.78 1024.0601 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1191.83 290.07 L1189.92 291.1 L1175.36 334.49 L1186.42 346.77 L1222.29 322.28 L1220.04 304.43 L1191.83 290.07 Z"
      /><path d="M1191.83 290.07 L1189.92 291.1 L1175.36 334.49 L1186.42 346.77 L1222.29 322.28 L1220.04 304.43 L1191.83 290.07 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1470.66 552.84 L1443.35 534.39 L1432.27 537.64 L1418.15 562.85 L1447.5601 592.15 L1466.65 588.2 L1470.66 552.84 Z"
      /><path d="M1470.66 552.84 L1443.35 534.39 L1432.27 537.64 L1418.15 562.85 L1447.5601 592.15 L1466.65 588.2 L1470.66 552.84 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M0 312.9 L35.12 316.65 L41.21 346.68 L19.11 370.74 L0 370.1 L0 312.9 Z"
      /><path d="M0 312.9 L35.12 316.65 L41.21 346.68 L19.11 370.74 L0 370.1 L0 312.9 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M85.23 799.7 L99.61 809.61 L90.25 850.42 L51.24 843.16 L44.8 827.22 L58.08 801.99 L85.23 799.7 Z"
      /><path d="M85.23 799.7 L99.61 809.61 L90.25 850.42 L51.24 843.16 L44.8 827.22 L58.08 801.99 L85.23 799.7 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M790.08 158.31 L829.16 165.32 L829.87 167.12 L813.92 198.14 L780.35 187.15 L790.08 158.31 Z"
      /><path d="M790.08 158.31 L829.16 165.32 L829.87 167.12 L813.92 198.14 L780.35 187.15 L790.08 158.31 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M859.8 411.53 L874.91 434.17 L872.73 446.1 L840.16 473.4 L813.08 459.91 L812.22 414.83 L819.78 407.99 L859.8 411.53 Z"
      /><path d="M859.8 411.53 L874.91 434.17 L872.73 446.1 L840.16 473.4 L813.08 459.91 L812.22 414.83 L819.78 407.99 L859.8 411.53 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M643.93 158.54 L614.45 162.96 L606.38 186.7 L616.83 198.8 L649.11 195.35 L653.69 168.06 L643.93 158.54 Z"
      /><path d="M643.93 158.54 L614.45 162.96 L606.38 186.7 L616.83 198.8 L649.11 195.35 L653.69 168.06 L643.93 158.54 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1361.48 608.27 L1386.5699 630.94 L1370.24 666.27 L1334.5601 639.57 L1344.36 612.57 L1361.48 608.27 Z"
      /><path d="M1361.48 608.27 L1386.5699 630.94 L1370.24 666.27 L1334.5601 639.57 L1344.36 612.57 L1361.48 608.27 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1288.99 415.46 L1262.85 415.31 L1249.37 437.67 L1264.63 465.53 L1300.75 462.61 L1307.8199 451.9 L1288.99 415.46 Z"
      /><path d="M1288.99 415.46 L1262.85 415.31 L1249.37 437.67 L1264.63 465.53 L1300.75 462.61 L1307.8199 451.9 L1288.99 415.46 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1578.22 340.14 L1546.6801 316.56 L1523.41 320.71 L1530.04 358.66 L1560.0601 365.1 L1576.6801 351.18 L1578.22 340.14 Z"
      /><path d="M1578.22 340.14 L1546.6801 316.56 L1523.41 320.71 L1530.04 358.66 L1560.0601 365.1 L1576.6801 351.18 L1578.22 340.14 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1810.76 52.93 L1839.3101 70.88 L1821.16 109.76 L1807.24 111.73 L1789.02 73.93 L1810.76 52.93 Z"
      /><path d="M1810.76 52.93 L1839.3101 70.88 L1821.16 109.76 L1807.24 111.73 L1789.02 73.93 L1810.76 52.93 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1561.7 398.51 L1571.2 403.82 L1579.85 423.74 L1547.35 451.51 L1543.2 449.96 L1533.52 431.66 L1544.29 403.91 L1561.7 398.51 Z"
      /><path d="M1561.7 398.51 L1571.2 403.82 L1579.85 423.74 L1547.35 451.51 L1543.2 449.96 L1533.52 431.66 L1544.29 403.91 L1561.7 398.51 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M820.08 1029.89 L778.2 1016.46 L769.07 1026.8101 L775.5 1080 L818.2 1080 L820.08 1029.89 Z"
      /><path d="M820.08 1029.89 L778.2 1016.46 L769.07 1026.8101 L775.5 1080 L818.2 1080 L820.08 1029.89 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M358.19 1034.9 L288.96 1022.34 L280.93 1029.77 L278 1080 L358.6 1080 L358.19 1034.9 Z"
      /><path d="M358.19 1034.9 L288.96 1022.34 L280.93 1029.77 L278 1080 L358.6 1080 L358.19 1034.9 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M216.28 745.45 L218.83 756.49 L193.45 801.26 L173.24 794.54 L159.68 762.89 L192.91 741.55 L216.28 745.45 Z"
      /><path d="M216.28 745.45 L218.83 756.49 L193.45 801.26 L173.24 794.54 L159.68 762.89 L192.91 741.55 L216.28 745.45 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M747.88 278.67 L700.68 290.37 L698.14 295.6 L700.69 307.47 L733.03 329.54 L755.29 308.93 L747.88 278.67 Z"
      /><path d="M747.88 278.67 L700.68 290.37 L698.14 295.6 L700.69 307.47 L733.03 329.54 L755.29 308.93 L747.88 278.67 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M69.73 751.45 L87.57 760.52 L85.23 799.7 L58.08 801.99 L44.32 779.36 L69.73 751.45 Z"
      /><path d="M69.73 751.45 L87.57 760.52 L85.23 799.7 L58.08 801.99 L44.32 779.36 L69.73 751.45 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M873.69 377.34 L859.8 411.53 L874.91 434.17 L913.56 420.96 L918.25 383.69 L916.58 381.47 L873.69 377.34 Z"
      /><path d="M873.69 377.34 L859.8 411.53 L874.91 434.17 L913.56 420.96 L918.25 383.69 L916.58 381.47 L873.69 377.34 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1355.6801 389.41 L1392.42 393.75 L1396.95 405.91 L1382.34 447.77 L1376.49 451.74 L1356.74 452.47 L1343.2 443.54 L1340.59 403.63 L1355.6801 389.41 Z"
      /><path d="M1355.6801 389.41 L1392.42 393.75 L1396.95 405.91 L1382.34 447.77 L1376.49 451.74 L1356.74 452.47 L1343.2 443.54 L1340.59 403.63 L1355.6801 389.41 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1148.63 538.72 L1115.49 543.31 L1115.96 588.32 L1152.26 586.65 L1160.59 548.29 L1148.63 538.72 Z"
      /><path d="M1148.63 538.72 L1115.49 543.31 L1115.96 588.32 L1152.26 586.65 L1160.59 548.29 L1148.63 538.72 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1766.95 335.08 L1742.8 376.59 L1703.4399 332.07 L1703.45 330.84 L1723.52 308.33 L1739.86 308.22 L1766.95 335.08 Z"
      /><path d="M1766.95 335.08 L1742.8 376.59 L1703.4399 332.07 L1703.45 330.84 L1723.52 308.33 L1739.86 308.22 L1766.95 335.08 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1023.8 549.93 L1048.9301 574.04 L1044.1 592.7 L1004.55 613.8 L984.45 585.74 L1000.48 552.85 L1023.8 549.93 Z"
      /><path d="M1023.8 549.93 L1048.9301 574.04 L1044.1 592.7 L1004.55 613.8 L984.45 585.74 L1000.48 552.85 L1023.8 549.93 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1647.38 652.72 L1621.87 663.8 L1615.59 699.49 L1630.04 717.57 L1656.27 706.76 L1671.25 664.74 L1647.38 652.72 Z"
      /><path d="M1647.38 652.72 L1621.87 663.8 L1615.59 699.49 L1630.04 717.57 L1656.27 706.76 L1671.25 664.74 L1647.38 652.72 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M614.82 221.7 L634.3 237.31 L634.66 239.16 L622.21 261.34 L609.28 265.25 L587.95 243.66 L587.74 234.41 L614.82 221.7 Z"
      /><path d="M614.82 221.7 L634.3 237.31 L634.66 239.16 L622.21 261.34 L609.28 265.25 L587.95 243.66 L587.74 234.41 L614.82 221.7 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M848.07 737.57 L883.46 764.73 L879.6 777.64 L838.73 793.09 L825.18 781.71 L832.32 740.36 L848.07 737.57 Z"
      /><path d="M848.07 737.57 L883.46 764.73 L879.6 777.64 L838.73 793.09 L825.18 781.71 L832.32 740.36 L848.07 737.57 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1870.74 118.59 L1911.01 157.27 L1860.7 183.37 L1840.87 166.19 L1849.27 127.73 L1870.74 118.59 Z"
      /><path d="M1870.74 118.59 L1911.01 157.27 L1860.7 183.37 L1840.87 166.19 L1849.27 127.73 L1870.74 118.59 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1192.15 145.76 L1160.98 117.95 L1128.9399 134.34 L1129.22 162.93 L1143.4 177.01 L1192.65 164.59 L1192.15 145.76 Z"
      /><path d="M1192.15 145.76 L1160.98 117.95 L1128.9399 134.34 L1129.22 162.93 L1143.4 177.01 L1192.65 164.59 L1192.15 145.76 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M438.35 161.08 L456.13 184.28 L439.9 212.21 L402.33 197.04 L400.17 170.57 L416.78 159.49 L438.35 161.08 Z"
      /><path d="M438.35 161.08 L456.13 184.28 L439.9 212.21 L402.33 197.04 L400.17 170.57 L416.78 159.49 L438.35 161.08 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M175.47 444.2 L150.27 406.01 L123.88 412.87 L116.79 424.3 L133.07 464.99 L138.65 468.73 L145.36 468.54 L166.41 458.72 L175.38 445.92 L175.47 444.2 Z"
      /><path d="M175.47 444.2 L150.27 406.01 L123.88 412.87 L116.79 424.3 L133.07 464.99 L138.65 468.73 L145.36 468.54 L166.41 458.72 L175.38 445.92 L175.47 444.2 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M736.44 228.16 L709.84 216.41 L699.68 221.61 L699.26 253.72 L731.42 250.36 L736.44 228.16 Z"
      /><path d="M736.44 228.16 L709.84 216.41 L699.68 221.61 L699.26 253.72 L731.42 250.36 L736.44 228.16 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1270.79 364.93 L1299.5 369.69 L1306.09 395.11 L1288.99 415.46 L1262.85 415.31 L1250.6899 392.88 L1270.79 364.93 Z"
      /><path d="M1270.79 364.93 L1299.5 369.69 L1306.09 395.11 L1288.99 415.46 L1262.85 415.31 L1250.6899 392.88 L1270.79 364.93 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M736.25 598.88 L710.88 571.75 L695.36 575.01 L683.86 608.36 L701.91 621.12 L736.25 598.88 Z"
      /><path d="M736.25 598.88 L710.88 571.75 L695.36 575.01 L683.86 608.36 L701.91 621.12 L736.25 598.88 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M914.01 105.38 L897.16 101.89 L869.37 120.26 L867.53 127.88 L886.75 162.05 L901.98 163.58 L930.18 131.54 L914.01 105.38 Z"
      /><path d="M914.01 105.38 L897.16 101.89 L869.37 120.26 L867.53 127.88 L886.75 162.05 L901.98 163.58 L930.18 131.54 L914.01 105.38 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1562.77 202.96 L1595.8199 218.17 L1599.98 247.03 L1565.6899 268.2 L1557.05 263.13 L1547.48 220.29 L1562.77 202.96 Z"
      /><path d="M1562.77 202.96 L1595.8199 218.17 L1599.98 247.03 L1565.6899 268.2 L1557.05 263.13 L1547.48 220.29 L1562.77 202.96 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1122.62 263.84 L1106.86 291.26 L1097.03 295.61 L1065.58 283.38 L1066.9399 244.95 L1122.62 263.84 Z"
      /><path d="M1122.62 263.84 L1106.86 291.26 L1097.03 295.61 L1065.58 283.38 L1066.9399 244.95 L1122.62 263.84 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1609.1801 379.36 L1576.6801 351.18 L1560.0601 365.1 L1561.7 398.51 L1571.2 403.82 L1609.1801 379.36 Z"
      /><path d="M1609.1801 379.36 L1576.6801 351.18 L1560.0601 365.1 L1561.7 398.51 L1571.2 403.82 L1609.1801 379.36 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1800.54 395.43 L1747.1 385.24 L1737.37 425.31 L1757.6 447.79 L1790.8 447.52 L1800.54 395.43 Z"
      /><path d="M1800.54 395.43 L1747.1 385.24 L1737.37 425.31 L1757.6 447.79 L1790.8 447.52 L1800.54 395.43 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1559.1899 119.08 L1575.74 129.81 L1580.85 163.09 L1560.88 185.1 L1523.46 165.28 L1523.54 140.17 L1559.1899 119.08 Z"
      /><path d="M1559.1899 119.08 L1575.74 129.81 L1580.85 163.09 L1560.88 185.1 L1523.46 165.28 L1523.54 140.17 L1559.1899 119.08 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1462.87 928.99 L1437.28 933.22 L1424.26 970.19 L1464.26 992.39 L1486.05 973.14 L1462.87 928.99 Z"
      /><path d="M1462.87 928.99 L1437.28 933.22 L1424.26 970.19 L1464.26 992.39 L1486.05 973.14 L1462.87 928.99 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M716.54 737.73 L670.4 745.89 L668.55 764 L712.84 797.22 L720.96 795.79 L735.26 763.18 L716.54 737.73 Z"
      /><path d="M716.54 737.73 L670.4 745.89 L668.55 764 L712.84 797.22 L720.96 795.79 L735.26 763.18 L716.54 737.73 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M581.58 791.17 L559.85 801.51 L557.72 850.34 L587.79 853.63 L611.19 829.03 L581.58 791.17 Z"
      /><path d="M581.58 791.17 L559.85 801.51 L557.72 850.34 L587.79 853.63 L611.19 829.03 L581.58 791.17 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M864.67 209.5 L894.37 223.33 L894.81 254.37 L856.18 266.75 L848.98 261.93 L851.83 218.36 L864.67 209.5 Z"
      /><path d="M864.67 209.5 L894.37 223.33 L894.81 254.37 L856.18 266.75 L848.98 261.93 L851.83 218.36 L864.67 209.5 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M953.77 978.73 L960.66 981.97 L966.98 991.76 L958.73 1028.3101 L924.77 1034.8199 L920.4 1029.73 L921.12 989.13 L953.77 978.73 Z"
      /><path d="M953.77 978.73 L960.66 981.97 L966.98 991.76 L958.73 1028.3101 L924.77 1034.8199 L920.4 1029.73 L921.12 989.13 L953.77 978.73 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1498.96 797.5 L1482.1 828.76 L1486.12 842.94 L1513.28 854.83 L1545.12 818.14 L1536.91 803.11 L1498.96 797.5 Z"
      /><path d="M1498.96 797.5 L1482.1 828.76 L1486.12 842.94 L1513.28 854.83 L1545.12 818.14 L1536.91 803.11 L1498.96 797.5 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M550.84 594.4 L563.53 596.4 L571.75 636.2 L546.15 642.13 L529.66 623 L550.84 594.4 Z"
      /><path d="M550.84 594.4 L563.53 596.4 L571.75 636.2 L546.15 642.13 L529.66 623 L550.84 594.4 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1166.59 764.65 L1138.3 750.84 L1111.4301 775.43 L1136.13 809.13 L1143.8 810.8 L1171 775.25 L1166.59 764.65 Z"
      /><path d="M1166.59 764.65 L1138.3 750.84 L1111.4301 775.43 L1136.13 809.13 L1143.8 810.8 L1171 775.25 L1166.59 764.65 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1863.85 580.03 L1870.65 633.44 L1809.28 636.85 L1801.49 611.6 L1814.04 583.98 L1863.85 580.03 Z"
      /><path d="M1863.85 580.03 L1870.65 633.44 L1809.28 636.85 L1801.49 611.6 L1814.04 583.98 L1863.85 580.03 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M175.38 445.92 L166.41 458.72 L187.54 491.78 L214.8 486.24 L217.26 464.71 L175.38 445.92 Z"
      /><path d="M175.38 445.92 L166.41 458.72 L187.54 491.78 L214.8 486.24 L217.26 464.71 L175.38 445.92 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M508.77 895.99 L496.15 923.11 L440 896.48 L442.61 882.65 L487 855.96 L508.77 895.99 Z"
      /><path d="M508.77 895.99 L496.15 923.11 L440 896.48 L442.61 882.65 L487 855.96 L508.77 895.99 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1544.77 42.56 L1496.8 33.13 L1482.29 56.07 L1505.4301 86.27 L1538.33 79.6 L1544.77 42.56 Z"
      /><path d="M1544.77 42.56 L1496.8 33.13 L1482.29 56.07 L1505.4301 86.27 L1538.33 79.6 L1544.77 42.56 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M281.79 398.92 L274.21 418.89 L229.99 424.11 L216.17 408.5 L215.59 404.28 L236.45 382.13 L263.92 382.07 L281.79 398.92 Z"
      /><path d="M281.79 398.92 L274.21 418.89 L229.99 424.11 L216.17 408.5 L215.59 404.28 L236.45 382.13 L263.92 382.07 L281.79 398.92 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M594.41 126.09 L551.01 110.14 L530.38 131.69 L531.89 137.62 L566.1 159.18 L594.21 134.31 L595.02 127.31 L594.41 126.09 Z"
      /><path d="M594.41 126.09 L551.01 110.14 L530.38 131.69 L531.89 137.62 L566.1 159.18 L594.21 134.31 L595.02 127.31 L594.41 126.09 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1329.26 689.46 L1320.4399 710.4 L1285.9301 702.16 L1278.47 676.99 L1310.23 661.36 L1329.26 689.46 Z"
      /><path d="M1329.26 689.46 L1320.4399 710.4 L1285.9301 702.16 L1278.47 676.99 L1310.23 661.36 L1329.26 689.46 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M705.64 514.71 L706.84 524.28 L670.14 550.3 L653.06 533.78 L652.42 523.5 L678.31 499.37 L705.64 514.71 Z"
      /><path d="M705.64 514.71 L706.84 524.28 L670.14 550.3 L653.06 533.78 L652.42 523.5 L678.31 499.37 L705.64 514.71 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M622.21 261.34 L650.41 287.31 L650.55 288.65 L614.26 305.08 L602.07 282.65 L609.28 265.25 L622.21 261.34 Z"
      /><path d="M622.21 261.34 L650.41 287.31 L650.55 288.65 L614.26 305.08 L602.07 282.65 L609.28 265.25 L622.21 261.34 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M267.22 620.04 L280.97 629.96 L284.04 650.54 L254.45 675.29 L240.03 670.7 L228.11 632.16 L267.22 620.04 Z"
      /><path d="M267.22 620.04 L280.97 629.96 L284.04 650.54 L254.45 675.29 L240.03 670.7 L228.11 632.16 L267.22 620.04 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1530.04 358.66 L1560.0601 365.1 L1561.7 398.51 L1544.29 403.91 L1517.8 387.69 L1515.95 374.92 L1530.04 358.66 Z"
      /><path d="M1530.04 358.66 L1560.0601 365.1 L1561.7 398.51 L1544.29 403.91 L1517.8 387.69 L1515.95 374.92 L1530.04 358.66 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1043.62 789.99 L1074.79 807.8 L1077.47 818.44 L1051.78 847.65 L1024.46 838.68 L1018.94 822.52 L1043.62 789.99 Z"
      /><path d="M1043.62 789.99 L1074.79 807.8 L1077.47 818.44 L1051.78 847.65 L1024.46 838.68 L1018.94 822.52 L1043.62 789.99 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M439.12 360.82 L465.77 368.46 L472.55 390.49 L461.13 408.55 L441.66 412.86 L422.51 386.7 L439.12 360.82 Z"
      /><path d="M439.12 360.82 L465.77 368.46 L472.55 390.49 L461.13 408.55 L441.66 412.86 L422.51 386.7 L439.12 360.82 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M271.25 342.21 L263.92 382.07 L281.79 398.92 L288.51 396.82 L308.51 369.58 L301 346.71 L271.25 342.21 Z"
      /><path d="M271.25 342.21 L263.92 382.07 L281.79 398.92 L288.51 396.82 L308.51 369.58 L301 346.71 L271.25 342.21 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1001.96 440.1 L988.24 486.52 L1042.7 503.74 L1044.89 502.75 L1061.63 461.44 L1054.6 446.76 L1001.96 440.1 Z"
      /><path d="M1001.96 440.1 L988.24 486.52 L1042.7 503.74 L1044.89 502.75 L1061.63 461.44 L1054.6 446.76 L1001.96 440.1 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M37.9 731.92 L67.92 746.7 L69.73 751.45 L44.32 779.36 L36.14 777.41 L18.75 746.32 L37.9 731.92 Z"
      /><path d="M37.9 731.92 L67.92 746.7 L69.73 751.45 L44.32 779.36 L36.14 777.41 L18.75 746.32 L37.9 731.92 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M981.49 43.76 L966.81 77.92 L938.93 73.22 L925 49.55 L956.71 10.66 L981.49 43.76 Z"
      /><path d="M981.49 43.76 L966.81 77.92 L938.93 73.22 L925 49.55 L956.71 10.66 L981.49 43.76 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M665.33 33.02 L678.81 46.7 L679.61 72.31 L644.65 89.57 L626.47 76.3 L626.81 47.71 L665.33 33.02 Z"
      /><path d="M665.33 33.02 L678.81 46.7 L679.61 72.31 L644.65 89.57 L626.47 76.3 L626.81 47.71 L665.33 33.02 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M652.42 523.5 L632.24 506.24 L605.5 519.91 L605.73 532.69 L625.07 549.59 L653.06 533.78 L652.42 523.5 Z"
      /><path d="M652.42 523.5 L632.24 506.24 L605.5 519.91 L605.73 532.69 L625.07 549.59 L653.06 533.78 L652.42 523.5 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1297.61 144.82 L1305.84 156.58 L1299.5 175.74 L1259.36 186.73 L1247.72 167.9 L1254.64 141.09 L1297.61 144.82 Z"
      /><path d="M1297.61 144.82 L1305.84 156.58 L1299.5 175.74 L1259.36 186.73 L1247.72 167.9 L1254.64 141.09 L1297.61 144.82 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M295.06 983.73 L253.69 952.19 L245.17 954.12 L224.75 984.05 L227.84 1014.05 L280.93 1029.77 L288.96 1022.34 L295.06 983.73 Z"
      /><path d="M295.06 983.73 L253.69 952.19 L245.17 954.12 L224.75 984.05 L227.84 1014.05 L280.93 1029.77 L288.96 1022.34 L295.06 983.73 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M44.32 779.36 L36.14 777.41 L0 800.1 L0 816.6 L44.8 827.22 L58.08 801.99 L44.32 779.36 Z"
      /><path d="M44.32 779.36 L36.14 777.41 L0 800.1 L0 816.6 L44.8 827.22 L58.08 801.99 L44.32 779.36 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1320.4399 710.4 L1327.24 732.39 L1326.7 732.88 L1289.79 743.38 L1269.4 725.03 L1285.9301 702.16 L1320.4399 710.4 Z"
      /><path d="M1320.4399 710.4 L1327.24 732.39 L1326.7 732.88 L1289.79 743.38 L1269.4 725.03 L1285.9301 702.16 L1320.4399 710.4 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1384.1899 224 L1433.16 226.39 L1439.97 232.47 L1428.72 265.91 L1385.4301 280.58 L1383.7 280.18 L1381.8199 277.55 L1378.5601 229.68 L1384.1899 224 Z"
      /><path d="M1384.1899 224 L1433.16 226.39 L1439.97 232.47 L1428.72 265.91 L1385.4301 280.58 L1383.7 280.18 L1381.8199 277.55 L1378.5601 229.68 L1384.1899 224 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M818.62 653.73 L840.07 679.27 L813.9 707.14 L783.58 687.58 L787.13 665.4 L818.62 653.73 Z"
      /><path d="M818.62 653.73 L840.07 679.27 L813.9 707.14 L783.58 687.58 L787.13 665.4 L818.62 653.73 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M97.74 131.52 L85.82 81.08 L53.35 86.93 L40.4 117 L49.25 130.53 L97.36 132.02 L97.74 131.52 Z"
      /><path d="M97.74 131.52 L85.82 81.08 L53.35 86.93 L40.4 117 L49.25 130.53 L97.36 132.02 L97.74 131.52 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1067.77 922.53 L1041.86 895.96 L1020.96 927.31 L1030.2 946.16 L1041.51 949 L1067.77 922.53 Z"
      /><path d="M1067.77 922.53 L1041.86 895.96 L1020.96 927.31 L1030.2 946.16 L1041.51 949 L1067.77 922.53 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M606.38 186.7 L583.44 189.71 L574.27 221.62 L587.74 234.41 L614.82 221.7 L616.83 198.8 L606.38 186.7 Z"
      /><path d="M606.38 186.7 L583.44 189.71 L574.27 221.62 L587.74 234.41 L614.82 221.7 L616.83 198.8 L606.38 186.7 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1660.9301 101.88 L1624.17 70.68 L1614.66 71.38 L1607.83 117.67 L1637.29 139.33 L1649.3199 135.7 L1660.9301 101.88 Z"
      /><path d="M1660.9301 101.88 L1624.17 70.68 L1614.66 71.38 L1607.83 117.67 L1637.29 139.33 L1649.3199 135.7 L1660.9301 101.88 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1392.65 570.82 L1413.87 623.79 L1386.5699 630.94 L1361.48 608.27 L1378.96 569.67 L1381.9301 568.38 L1392.65 570.82 Z"
      /><path d="M1392.65 570.82 L1413.87 623.79 L1386.5699 630.94 L1361.48 608.27 L1378.96 569.67 L1381.9301 568.38 L1392.65 570.82 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1179.35 992.63 L1213.87 1013.05 L1217.1801 1030.77 L1179 1048.79 L1168.14 1038.9301 L1179.35 992.63 Z"
      /><path d="M1179.35 992.63 L1213.87 1013.05 L1217.1801 1030.77 L1179 1048.79 L1168.14 1038.9301 L1179.35 992.63 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M902.53 961.55 L864.75 950.28 L851.48 1006.7 L852.39 1009.18 L856.7 1011.05 L905.6 976.68 L902.53 961.55 Z"
      /><path d="M902.53 961.55 L864.75 950.28 L851.48 1006.7 L852.39 1009.18 L856.7 1011.05 L905.6 976.68 L902.53 961.55 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M133.07 464.99 L116.79 424.3 L85.3 433.9 L84.67 467.94 L91.3 472.64 L133.07 464.99 Z"
      /><path d="M133.07 464.99 L116.79 424.3 L85.3 433.9 L84.67 467.94 L91.3 472.64 L133.07 464.99 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M256.9 41.73 L274.97 56.33 L274.35 79.86 L239.96 106.08 L238.02 106.29 L228.9 100.96 L221.2 55.86 L256.9 41.73 Z"
      /><path d="M256.9 41.73 L274.97 56.33 L274.35 79.86 L239.96 106.08 L238.02 106.29 L228.9 100.96 L221.2 55.86 L256.9 41.73 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1038.02 994.45 L1045.24 1030.39 L1037.62 1037.02 L1002.39 1031.47 L1001.39 996.75 L1010.54 988.64 L1038.02 994.45 Z"
      /><path d="M1038.02 994.45 L1045.24 1030.39 L1037.62 1037.02 L1002.39 1031.47 L1001.39 996.75 L1010.54 988.64 L1038.02 994.45 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M146.04 44.13 L101.48 32.57 L89.62 45.36 L90.17 75.96 L133.46 81.79 L153.48 60.47 L146.04 44.13 Z"
      /><path d="M146.04 44.13 L101.48 32.57 L89.62 45.36 L90.17 75.96 L133.46 81.79 L153.48 60.47 L146.04 44.13 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M656.1 330.73 L635.26 337.81 L623.43 366.86 L627.61 378.97 L673.8 376.15 L679.89 348.47 L677.02 341.68 L656.1 330.73 Z"
      /><path d="M656.1 330.73 L635.26 337.81 L623.43 366.86 L627.61 378.97 L673.8 376.15 L679.89 348.47 L677.02 341.68 L656.1 330.73 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M541 489.5 L541.1 512.38 L522.64 523.84 L490.63 511.49 L490.43 502.02 L509.55 477.17 L523.72 474.55 L541 489.5 Z"
      /><path d="M541 489.5 L541.1 512.38 L522.64 523.84 L490.63 511.49 L490.43 502.02 L509.55 477.17 L523.72 474.55 L541 489.5 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M808.99 29.99 L844.4 41.76 L845.28 54.12 L809.08 71.91 L793.01 61.65 L790.42 45.49 L808.99 29.99 Z"
      /><path d="M808.99 29.99 L844.4 41.76 L845.28 54.12 L809.08 71.91 L793.01 61.65 L790.42 45.49 L808.99 29.99 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M522.95 305.37 L484.25 299.79 L469.37 317.29 L487.76 345.7 L492.28 346.4 L516.77 333.37 L524.92 308.38 L522.95 305.37 Z"
      /><path d="M522.95 305.37 L484.25 299.79 L469.37 317.29 L487.76 345.7 L492.28 346.4 L516.77 333.37 L524.92 308.38 L522.95 305.37 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1126.7 678.55 L1093.29 670.76 L1089.38 673.18 L1080.78 714.46 L1087.5699 723.77 L1127.3199 720.01 L1126.7 678.55 Z"
      /><path d="M1126.7 678.55 L1093.29 670.76 L1089.38 673.18 L1080.78 714.46 L1087.5699 723.77 L1127.3199 720.01 L1126.7 678.55 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M679.89 348.47 L673.8 376.15 L681.7 388.01 L720 385.76 L733.23 356.72 L731.27 352.79 L679.89 348.47 Z"
      /><path d="M679.89 348.47 L673.8 376.15 L681.7 388.01 L720 385.76 L733.23 356.72 L731.27 352.79 L679.89 348.47 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1513.97 707.88 L1477.71 727.07 L1498.38 760.99 L1531.23 751.05 L1535.12 737.48 L1513.97 707.88 Z"
      /><path d="M1513.97 707.88 L1477.71 727.07 L1498.38 760.99 L1531.23 751.05 L1535.12 737.48 L1513.97 707.88 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1839.22 8.9 L1856.4 28.65 L1853.9399 68.19 L1839.3101 70.88 L1810.76 52.93 L1809.65 43.62 L1839.22 8.9 Z"
      /><path d="M1839.22 8.9 L1856.4 28.65 L1853.9399 68.19 L1839.3101 70.88 L1810.76 52.93 L1809.65 43.62 L1839.22 8.9 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1089.84 179.95 L1090.9399 208.97 L1065.25 231.04 L1034.0699 196.01 L1056.55 162.49 L1064.64 160.66 L1089.84 179.95 Z"
      /><path d="M1089.84 179.95 L1090.9399 208.97 L1065.25 231.04 L1034.0699 196.01 L1056.55 162.49 L1064.64 160.66 L1089.84 179.95 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1920 565 L1920 494.1 L1858.72 507.52 L1852.28 518.53 L1873.28 568.3 L1920 565 Z"
      /><path d="M1920 565 L1920 494.1 L1858.72 507.52 L1852.28 518.53 L1873.28 568.3 L1920 565 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1894.2 56.21 L1920 70.5 L1920 85.1 L1875.45 105.09 L1856.04 69.2 L1894.2 56.21 Z"
      /><path d="M1894.2 56.21 L1920 70.5 L1920 85.1 L1875.45 105.09 L1856.04 69.2 L1894.2 56.21 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1680.6 807.24 L1670.9301 823.76 L1635.51 834.15 L1628.54 831.63 L1621.48 788.64 L1646.51 772.51 L1680.6 807.24 Z"
      /><path d="M1680.6 807.24 L1670.9301 823.76 L1635.51 834.15 L1628.54 831.63 L1621.48 788.64 L1646.51 772.51 L1680.6 807.24 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1806.24 225.52 L1821.25 232.97 L1825.05 279.94 L1797.85 290.99 L1767.45 272.3 L1761.73 252.06 L1806.24 225.52 Z"
      /><path d="M1806.24 225.52 L1821.25 232.97 L1825.05 279.94 L1797.85 290.99 L1767.45 272.3 L1761.73 252.06 L1806.24 225.52 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M487.76 345.7 L465.77 368.46 L472.55 390.49 L511.38 393.32 L514.05 381.91 L492.28 346.4 L487.76 345.7 Z"
      /><path d="M487.76 345.7 L465.77 368.46 L472.55 390.49 L511.38 393.32 L514.05 381.91 L492.28 346.4 L487.76 345.7 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M983.47 939.39 L968.14 934.33 L945.05 944.77 L953.77 978.73 L960.66 981.97 L988.39 954.11 L983.47 939.39 Z"
      /><path d="M983.47 939.39 L968.14 934.33 L945.05 944.77 L953.77 978.73 L960.66 981.97 L988.39 954.11 L983.47 939.39 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M51.24 843.16 L34.29 872.34 L56.19 900.29 L78.39 895.87 L95.87 858.52 L90.25 850.42 L51.24 843.16 Z"
      /><path d="M51.24 843.16 L34.29 872.34 L56.19 900.29 L78.39 895.87 L95.87 858.52 L90.25 850.42 L51.24 843.16 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M213.7 1080 L204.91 1039.0601 L145.1 1053.28 L141.2 1080 L213.7 1080 Z"
      /><path d="M213.7 1080 L204.91 1039.0601 L145.1 1053.28 L141.2 1080 L213.7 1080 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M20.62 483.83 L0 481.3 L0 537.1 L0.92 537.07 L35.48 513.66 L20.62 483.83 Z"
      /><path d="M20.62 483.83 L0 481.3 L0 537.1 L0.92 537.07 L35.48 513.66 L20.62 483.83 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1804.1 649.95 L1841.14 696.19 L1812.29 724.29 L1785.01 718.38 L1779.63 665.45 L1804.1 649.95 Z"
      /><path d="M1804.1 649.95 L1841.14 696.19 L1812.29 724.29 L1785.01 718.38 L1779.63 665.45 L1804.1 649.95 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M154.41 996.65 L135.54 1032.78 L99.7 1027.76 L91.49 995.71 L107.3 976.57 L154.41 996.65 Z"
      /><path d="M154.41 996.65 L135.54 1032.78 L99.7 1027.76 L91.49 995.71 L107.3 976.57 L154.41 996.65 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M383.11 302.43 L406.71 337.52 L387.03 356.63 L358.13 347.46 L374.39 301.88 L383.11 302.43 Z"
      /><path d="M383.11 302.43 L406.71 337.52 L387.03 356.63 L358.13 347.46 L374.39 301.88 L383.11 302.43 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M894.65 590.01 L905.57 599.27 L892.96 645.49 L877.51 649.41 L845.64 618.62 L852.86 597.26 L894.65 590.01 Z"
      /><path d="M894.65 590.01 L905.57 599.27 L892.96 645.49 L877.51 649.41 L845.64 618.62 L852.86 597.26 L894.65 590.01 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M41.21 346.68 L19.11 370.74 L37.52 390.99 L68.52 391.71 L89.08 368.52 L80.09 355 L41.21 346.68 Z"
      /><path d="M41.21 346.68 L19.11 370.74 L37.52 390.99 L68.52 391.71 L89.08 368.52 L80.09 355 L41.21 346.68 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M155.57 693.74 L128.51 698.36 L121.15 728.44 L144.66 735.18 L168.41 703.39 L155.57 693.74 Z"
      /><path d="M155.57 693.74 L128.51 698.36 L121.15 728.44 L144.66 735.18 L168.41 703.39 L155.57 693.74 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1396.9399 505.85 L1396.39 505.84 L1380.6899 515.7 L1381.9301 568.38 L1392.65 570.82 L1418.15 562.85 L1432.27 537.64 L1396.9399 505.85 Z"
      /><path d="M1396.9399 505.85 L1396.39 505.84 L1380.6899 515.7 L1381.9301 568.38 L1392.65 570.82 L1418.15 562.85 L1432.27 537.64 L1396.9399 505.85 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M561.23 907.15 L544.18 887.72 L508.77 895.99 L496.15 923.11 L496.32 923.97 L515.88 941.16 L556.12 931.42 L561.23 907.15 Z"
      /><path d="M561.23 907.15 L544.18 887.72 L508.77 895.99 L496.15 923.11 L496.32 923.97 L515.88 941.16 L556.12 931.42 L561.23 907.15 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1170.8 0 L1110.2 0 L1129.74 61.72 L1137.3199 62.67 L1173.0699 35.97 L1170.8 0 Z"
      /><path d="M1170.8 0 L1110.2 0 L1129.74 61.72 L1137.3199 62.67 L1173.0699 35.97 L1170.8 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M490.63 511.49 L522.64 523.84 L522.54 560.83 L483.64 555.68 L480.66 522.49 L490.63 511.49 Z"
      /><path d="M490.63 511.49 L522.64 523.84 L522.54 560.83 L483.64 555.68 L480.66 522.49 L490.63 511.49 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M713.58 85.72 L734.9 109.46 L733.39 121.2 L717.84 134.97 L686.77 127.14 L685.56 125.49 L696.63 87.05 L713.58 85.72 Z"
      /><path d="M713.58 85.72 L734.9 109.46 L733.39 121.2 L717.84 134.97 L686.77 127.14 L685.56 125.49 L696.63 87.05 L713.58 85.72 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M842.5 934.86 L807.29 963.98 L800.46 963.87 L781.72 937.38 L792.56 901.89 L826.23 901.28 L842.5 934.86 Z"
      /><path d="M842.5 934.86 L807.29 963.98 L800.46 963.87 L781.72 937.38 L792.56 901.89 L826.23 901.28 L842.5 934.86 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M475.22 747.21 L514.52 768.4 L515.71 781.42 L460.19 811.18 L455.38 809.48 L441.63 778.47 L475.22 747.21 Z"
      /><path d="M475.22 747.21 L514.52 768.4 L515.71 781.42 L460.19 811.18 L455.38 809.48 L441.63 778.47 L475.22 747.21 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M556.73 695.47 L536.49 724.49 L537.58 738.54 L593.53 760.72 L604.66 738.71 L602.21 715.47 L556.73 695.47 Z"
      /><path d="M556.73 695.47 L536.49 724.49 L537.58 738.54 L593.53 760.72 L604.66 738.71 L602.21 715.47 L556.73 695.47 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M953.81 877.1 L925.76 866.67 L916.75 886.74 L925.65 907.48 L934.54 910.42 L960.68 898.79 L953.81 877.1 Z"
      /><path d="M953.81 877.1 L925.76 866.67 L916.75 886.74 L925.65 907.48 L934.54 910.42 L960.68 898.79 L953.81 877.1 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M44.4 0 L0 0 L0 59.6 L30.34 58.6 L50.16 32.6 L44.4 0 Z"
      /><path d="M44.4 0 L0 0 L0 59.6 L30.34 58.6 L50.16 32.6 L44.4 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1632.8199 605.32 L1610.71 565.86 L1592.5 568.56 L1569.71 597.76 L1590.83 626.53 L1632.8199 605.32 Z"
      /><path d="M1632.8199 605.32 L1610.71 565.86 L1592.5 568.56 L1569.71 597.76 L1590.83 626.53 L1632.8199 605.32 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M869.37 120.26 L847.11 96.01 L816.09 102.58 L814.17 105.57 L815.31 122.68 L833.67 142.6 L867.53 127.88 L869.37 120.26 Z"
      /><path d="M869.37 120.26 L847.11 96.01 L816.09 102.58 L814.17 105.57 L815.31 122.68 L833.67 142.6 L867.53 127.88 L869.37 120.26 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1752.36 119.35 L1713.0601 101.7 L1708.21 102.79 L1693.27 155.34 L1721.6 164.96 L1748.7 144.97 L1752.36 119.35 Z"
      /><path d="M1752.36 119.35 L1713.0601 101.7 L1708.21 102.79 L1693.27 155.34 L1721.6 164.96 L1748.7 144.97 L1752.36 119.35 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1872.36 751.89 L1855.74 766.8 L1867.73 802.62 L1920 799 L1920 759.3 L1872.36 751.89 Z"
      /><path d="M1872.36 751.89 L1855.74 766.8 L1867.73 802.62 L1920 799 L1920 759.3 L1872.36 751.89 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1262.95 996.09 L1305.46 1006.07 L1297.21 1038.64 L1295.29 1039.72 L1260.28 1022.35 L1262.95 996.09 Z"
      /><path d="M1262.95 996.09 L1305.46 1006.07 L1297.21 1038.64 L1295.29 1039.72 L1260.28 1022.35 L1262.95 996.09 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M288.51 396.82 L281.79 398.92 L274.21 418.89 L280.83 439.21 L313.5 448.11 L332.83 426.99 L331.64 418.05 L288.51 396.82 Z"
      /><path d="M288.51 396.82 L281.79 398.92 L274.21 418.89 L280.83 439.21 L313.5 448.11 L332.83 426.99 L331.64 418.05 L288.51 396.82 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1386.0699 868.1 L1426.4399 872.21 L1418.38 916.55 L1385.63 920.86 L1372.73 903.18 L1386.0699 868.1 Z"
      /><path d="M1386.0699 868.1 L1426.4399 872.21 L1418.38 916.55 L1385.63 920.86 L1372.73 903.18 L1386.0699 868.1 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1797.85 290.99 L1767.45 272.3 L1739.86 308.22 L1766.95 335.08 L1790.3101 331.65 L1797.85 290.99 Z"
      /><path d="M1797.85 290.99 L1767.45 272.3 L1739.86 308.22 L1766.95 335.08 L1790.3101 331.65 L1797.85 290.99 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1391.6 774.3 L1391.86 774.86 L1380.27 823.74 L1379.0601 824.62 L1346.76 812.98 L1340.03 790.17 L1356 772.05 L1391.6 774.3 Z"
      /><path d="M1391.6 774.3 L1391.86 774.86 L1380.27 823.74 L1379.0601 824.62 L1346.76 812.98 L1340.03 790.17 L1356 772.05 L1391.6 774.3 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M85.62 663.37 L75.16 664.69 L73.37 704.49 L81.73 712.01 L87.33 711.81 L112.05 684.53 L111.16 679.68 L85.62 663.37 Z"
      /><path d="M85.62 663.37 L75.16 664.69 L73.37 704.49 L81.73 712.01 L87.33 711.81 L112.05 684.53 L111.16 679.68 L85.62 663.37 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1120.85 998.52 L1135.29 1002.51 L1147.22 1037.3199 L1128.62 1051.97 L1102.59 1034.1899 L1120.85 998.52 Z"
      /><path d="M1120.85 998.52 L1135.29 1002.51 L1147.22 1037.3199 L1128.62 1051.97 L1102.59 1034.1899 L1120.85 998.52 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1789.36 995.88 L1737.09 990.94 L1728.53 1004.45 L1731.23 1027.51 L1770.08 1043.25 L1788.9399 1026.83 L1789.36 995.88 Z"
      /><path d="M1789.36 995.88 L1737.09 990.94 L1728.53 1004.45 L1731.23 1027.51 L1770.08 1043.25 L1788.9399 1026.83 L1789.36 995.88 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1757.6 447.79 L1737.37 425.31 L1705.85 432.99 L1696.63 450.35 L1720.85 493.59 L1734.78 491.62 L1757.6 447.79 Z"
      /><path d="M1757.6 447.79 L1737.37 425.31 L1705.85 432.99 L1696.63 450.35 L1720.85 493.59 L1734.78 491.62 L1757.6 447.79 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M879.6 777.64 L894.66 809.32 L880.93 828.16 L841.43 814.2 L838.73 793.09 L879.6 777.64 Z"
      /><path d="M879.6 777.64 L894.66 809.32 L880.93 828.16 L841.43 814.2 L838.73 793.09 L879.6 777.64 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1803.25 393.57 L1835.27 398.19 L1857.52 440.85 L1842.1899 459.25 L1802.42 459.56 L1790.8 447.52 L1800.54 395.43 L1803.25 393.57 Z"
      /><path d="M1803.25 393.57 L1835.27 398.19 L1857.52 440.85 L1842.1899 459.25 L1802.42 459.56 L1790.8 447.52 L1800.54 395.43 L1803.25 393.57 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M783.82 144.85 L790.08 158.31 L780.35 187.15 L778.92 187.9 L750.89 180.08 L746.88 165.35 L763.11 141.46 L772.63 139.14 L783.82 144.85 Z"
      /><path d="M783.82 144.85 L790.08 158.31 L780.35 187.15 L778.92 187.9 L750.89 180.08 L746.88 165.35 L763.11 141.46 L772.63 139.14 L783.82 144.85 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M154.7 525.13 L126.08 499.72 L114.41 504.9 L112.73 529.84 L125.66 538.84 L154.7 525.13 Z"
      /><path d="M154.7 525.13 L126.08 499.72 L114.41 504.9 L112.73 529.84 L125.66 538.84 L154.7 525.13 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1042.7 503.74 L1023.8 549.93 L1000.48 552.85 L972.75 524.19 L979.39 491.81 L988.24 486.52 L1042.7 503.74 Z"
      /><path d="M1042.7 503.74 L1023.8 549.93 L1000.48 552.85 L972.75 524.19 L979.39 491.81 L988.24 486.52 L1042.7 503.74 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1317.04 839.46 L1315.73 838.9 L1274.61 849.34 L1268.97 868.47 L1283.85 894.29 L1328.86 865.23 L1317.04 839.46 Z"
      /><path d="M1317.04 839.46 L1315.73 838.9 L1274.61 849.34 L1268.97 868.47 L1283.85 894.29 L1328.86 865.23 L1317.04 839.46 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M740.8 191.59 L715.04 191.51 L709.84 216.41 L736.44 228.16 L745.46 222.01 L740.8 191.59 Z"
      /><path d="M740.8 191.59 L715.04 191.51 L709.84 216.41 L736.44 228.16 L745.46 222.01 L740.8 191.59 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1567.24 723.3 L1589.4399 748.92 L1586.36 768.71 L1547.01 774.53 L1531.23 751.05 L1535.12 737.48 L1567.24 723.3 Z"
      /><path d="M1567.24 723.3 L1589.4399 748.92 L1586.36 768.71 L1547.01 774.53 L1531.23 751.05 L1535.12 737.48 L1567.24 723.3 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M668.55 764 L712.84 797.22 L684.67 826.87 L647.05 797.98 L646.99 788.19 L668.55 764 Z"
      /><path d="M668.55 764 L712.84 797.22 L684.67 826.87 L647.05 797.98 L646.99 788.19 L668.55 764 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1256.41 55.33 L1259.03 66.54 L1222.41 100.04 L1200.3101 83.52 L1200.78 52.4 L1228.26 37.17 L1256.41 55.33 Z"
      /><path d="M1256.41 55.33 L1259.03 66.54 L1222.41 100.04 L1200.3101 83.52 L1200.78 52.4 L1228.26 37.17 L1256.41 55.33 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M480.66 522.49 L483.64 555.68 L465.9 574.22 L433.19 549.52 L433.22 528.29 L440.27 520.9 L480.66 522.49 Z"
      /><path d="M480.66 522.49 L483.64 555.68 L465.9 574.22 L433.19 549.52 L433.22 528.29 L440.27 520.9 L480.66 522.49 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1022.73 251.74 L998.56 227.28 L967.55 245.97 L981.05 283.61 L1016.47 280.2 L1022.73 251.74 Z"
      /><path d="M1022.73 251.74 L998.56 227.28 L967.55 245.97 L981.05 283.61 L1016.47 280.2 L1022.73 251.74 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1187.77 356.58 L1220.09 372.22 L1225.61 386.41 L1201.66 415.02 L1185.5699 413.55 L1166.71 383.8 L1187.77 356.58 Z"
      /><path d="M1187.77 356.58 L1220.09 372.22 L1225.61 386.41 L1201.66 415.02 L1185.5699 413.55 L1166.71 383.8 L1187.77 356.58 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M50.16 32.6 L30.34 58.6 L53.35 86.93 L85.82 81.08 L90.17 75.96 L89.62 45.36 L50.16 32.6 Z"
      /><path d="M50.16 32.6 L30.34 58.6 L53.35 86.93 L85.82 81.08 L90.17 75.96 L89.62 45.36 L50.16 32.6 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1446.8199 693.29 L1418.3101 716.35 L1379.4399 685.11 L1379.4301 685.07 L1428.92 662.82 L1446.8199 693.29 Z"
      /><path d="M1446.8199 693.29 L1418.3101 716.35 L1379.4399 685.11 L1379.4301 685.07 L1428.92 662.82 L1446.8199 693.29 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M166.41 458.72 L187.54 491.78 L175.66 513.11 L166.66 515.86 L145.36 468.54 L166.41 458.72 Z"
      /><path d="M166.41 458.72 L187.54 491.78 L175.66 513.11 L166.66 515.86 L145.36 468.54 L166.41 458.72 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M529.66 623 L501.58 621.08 L497 628.24 L508.44 668.63 L536.57 668.57 L546.15 642.13 L529.66 623 Z"
      /><path d="M529.66 623 L501.58 621.08 L497 628.24 L508.44 668.63 L536.57 668.57 L546.15 642.13 L529.66 623 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M123.87 565.17 L129.31 572.72 L118.5 594.74 L95.85 599.58 L79.98 581.27 L84 564.03 L90.45 560.05 L123.87 565.17 Z"
      /><path d="M123.87 565.17 L129.31 572.72 L118.5 594.74 L95.85 599.58 L79.98 581.27 L84 564.03 L90.45 560.05 L123.87 565.17 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M403.41 58.07 L415.43 64.45 L418.48 107.99 L410.23 114.44 L380.48 116.2 L374.04 110.31 L371 73.63 L379.28 61.24 L403.41 58.07 Z"
      /><path d="M403.41 58.07 L415.43 64.45 L418.48 107.99 L410.23 114.44 L380.48 116.2 L374.04 110.31 L371 73.63 L379.28 61.24 L403.41 58.07 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1643.22 201.78 L1627.9399 194.15 L1595.8199 218.17 L1599.98 247.03 L1624.54 259.1 L1644.85 246.27 L1643.22 201.78 Z"
      /><path d="M1643.22 201.78 L1627.9399 194.15 L1595.8199 218.17 L1599.98 247.03 L1624.54 259.1 L1644.85 246.27 L1643.22 201.78 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M323.42 784.99 L322.74 801.23 L287.2 816.13 L262.44 785.3 L284.39 757.45 L286.21 757.11 L323.42 784.99 Z"
      /><path d="M323.42 784.99 L322.74 801.23 L287.2 816.13 L262.44 785.3 L284.39 757.45 L286.21 757.11 L323.42 784.99 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M730.05 487.62 L705.64 514.71 L706.84 524.28 L723.43 543.07 L746.84 543.03 L769.17 513.28 L730.05 487.62 Z"
      /><path d="M730.05 487.62 L705.64 514.71 L706.84 524.28 L723.43 543.07 L746.84 543.03 L769.17 513.28 L730.05 487.62 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1043.42 652.95 L1044.83 662.1 L1033.46 678.97 L986.05 677.94 L981.35 644.98 L1003.36 623.23 L1043.42 652.95 Z"
      /><path d="M1043.42 652.95 L1044.83 662.1 L1033.46 678.97 L986.05 677.94 L981.35 644.98 L1003.36 623.23 L1043.42 652.95 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1885.53 941.28 L1861.58 905.02 L1825.4 934.44 L1839.33 961.89 L1871.77 962.79 L1885.53 941.28 Z"
      /><path d="M1885.53 941.28 L1861.58 905.02 L1825.4 934.44 L1839.33 961.89 L1871.77 962.79 L1885.53 941.28 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M601.86 1034.64 L590.03 996.39 L548.42 1006.69 L544.19 1022.5 L565.52 1046.7 L601.86 1034.64 Z"
      /><path d="M601.86 1034.64 L590.03 996.39 L548.42 1006.69 L544.19 1022.5 L565.52 1046.7 L601.86 1034.64 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M820.75 264.69 L806.92 279.76 L771.09 263.35 L776.4 231.33 L807.56 229.46 L820.75 264.69 Z"
      /><path d="M820.75 264.69 L806.92 279.76 L771.09 263.35 L776.4 231.33 L807.56 229.46 L820.75 264.69 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1024.6 0 L956.5 0 L956.71 10.66 L981.49 43.76 L1019.25 40.41 L1024.6 0 Z"
      /><path d="M1024.6 0 L956.5 0 L956.71 10.66 L981.49 43.76 L1019.25 40.41 L1024.6 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M659.57 209.16 L671.67 212.56 L669.94 254.08 L665.99 255.76 L634.66 239.16 L634.3 237.31 L659.57 209.16 Z"
      /><path d="M659.57 209.16 L671.67 212.56 L669.94 254.08 L665.99 255.76 L634.66 239.16 L634.3 237.31 L659.57 209.16 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1222.29 322.28 L1186.42 346.77 L1187.77 356.58 L1220.09 372.22 L1240.74 339.55 L1222.29 322.28 Z"
      /><path d="M1222.29 322.28 L1186.42 346.77 L1187.77 356.58 L1220.09 372.22 L1240.74 339.55 L1222.29 322.28 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M650.15 961.81 L678.49 962.32 L683.13 990.41 L670.24 1004.04 L635.2 989.26 L650.15 961.81 Z"
      /><path d="M650.15 961.81 L678.49 962.32 L683.13 990.41 L670.24 1004.04 L635.2 989.26 L650.15 961.81 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M133.07 464.99 L138.65 468.73 L126.08 499.72 L114.41 504.9 L97.23 497.89 L91.3 472.64 L133.07 464.99 Z"
      /><path d="M133.07 464.99 L138.65 468.73 L126.08 499.72 L114.41 504.9 L97.23 497.89 L91.3 472.64 L133.07 464.99 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1557.05 263.13 L1526.48 269.61 L1501.17 245.07 L1513.15 221 L1547.48 220.29 L1557.05 263.13 Z"
      /><path d="M1557.05 263.13 L1526.48 269.61 L1501.17 245.07 L1513.15 221 L1547.48 220.29 L1557.05 263.13 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1149.9 495.53 L1115.64 488.17 L1093.9399 527.93 L1115.49 543.31 L1148.63 538.72 L1149.9 495.53 Z"
      /><path d="M1149.9 495.53 L1115.64 488.17 L1093.9399 527.93 L1115.49 543.31 L1148.63 538.72 L1149.9 495.53 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M760.99 451.67 L789.84 469.84 L778.44 511.21 L769.17 513.28 L730.05 487.62 L728.78 472.97 L760.99 451.67 Z"
      /><path d="M760.99 451.67 L789.84 469.84 L778.44 511.21 L769.17 513.28 L730.05 487.62 L728.78 472.97 L760.99 451.67 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1477.71 727.07 L1474.9 726.32 L1445.17 750.44 L1450.5601 777.54 L1490.79 779.05 L1498.38 760.99 L1477.71 727.07 Z"
      /><path d="M1477.71 727.07 L1474.9 726.32 L1445.17 750.44 L1450.5601 777.54 L1490.79 779.05 L1498.38 760.99 L1477.71 727.07 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M306.12 488.08 L301.9 507.45 L276.79 517.99 L253.38 498.8 L265.48 471.98 L306.12 488.08 Z"
      /><path d="M306.12 488.08 L301.9 507.45 L276.79 517.99 L253.38 498.8 L265.48 471.98 L306.12 488.08 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1809.65 43.62 L1773.5601 18.05 L1750.5 54.93 L1767.3199 72.9 L1789.02 73.93 L1810.76 52.93 L1809.65 43.62 Z"
      /><path d="M1809.65 43.62 L1773.5601 18.05 L1750.5 54.93 L1767.3199 72.9 L1789.02 73.93 L1810.76 52.93 L1809.65 43.62 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1648.9 0 L1712.4 0 L1711.63 36.59 L1681.79 52.45 L1657.64 42.17 L1648.9 0 Z"
      /><path d="M1648.9 0 L1712.4 0 L1711.63 36.59 L1681.79 52.45 L1657.64 42.17 L1648.9 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M352.01 635.46 L342.26 634.64 L306.74 662.91 L315.31 692.92 L343.81 691.25 L356.94 648.7 L352.01 635.46 Z"
      /><path d="M352.01 635.46 L342.26 634.64 L306.74 662.91 L315.31 692.92 L343.81 691.25 L356.94 648.7 L352.01 635.46 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1083.6 0 L1110.2 0 L1129.74 61.72 L1112.25 72.32 L1070.41 63.91 L1066.78 58.68 L1083.6 0 Z"
      /><path d="M1083.6 0 L1110.2 0 L1129.74 61.72 L1112.25 72.32 L1070.41 63.91 L1066.78 58.68 L1083.6 0 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1017.44 136.34 L1056.55 162.49 L1034.0699 196.01 L1003.76 199.86 L999.01 194.34 L1001.79 146.38 L1017.44 136.34 Z"
      /><path d="M1017.44 136.34 L1056.55 162.49 L1034.0699 196.01 L1003.76 199.86 L999.01 194.34 L1001.79 146.38 L1017.44 136.34 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1598.03 52.39 L1550.71 37.38 L1544.77 42.56 L1538.33 79.6 L1555.86 96.13 L1604.86 65.37 L1598.03 52.39 Z"
      /><path d="M1598.03 52.39 L1550.71 37.38 L1544.77 42.56 L1538.33 79.6 L1555.86 96.13 L1604.86 65.37 L1598.03 52.39 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1761.73 252.06 L1749.1801 244.76 L1705.15 270.66 L1723.52 308.33 L1739.86 308.22 L1767.45 272.3 L1761.73 252.06 Z"
      /><path d="M1761.73 252.06 L1749.1801 244.76 L1705.15 270.66 L1723.52 308.33 L1739.86 308.22 L1767.45 272.3 L1761.73 252.06 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M560.9 0 L610.9 0 L609.89 33.14 L578.64 45.89 L562.5 33.46 L560.9 0 Z"
      /><path d="M560.9 0 L610.9 0 L609.89 33.14 L578.64 45.89 L562.5 33.46 L560.9 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M856.18 266.75 L848.98 261.93 L820.75 264.69 L806.92 279.76 L806.88 300.97 L836.76 318.2 L862.79 302.24 L856.18 266.75 Z"
      /><path d="M856.18 266.75 L848.98 261.93 L820.75 264.69 L806.92 279.76 L806.88 300.97 L836.76 318.2 L862.79 302.24 L856.18 266.75 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1228.9 0 L1284 0 L1286.88 22.57 L1256.41 55.33 L1228.26 37.17 L1228.9 0 Z"
      /><path d="M1228.9 0 L1284 0 L1286.88 22.57 L1256.41 55.33 L1228.26 37.17 L1228.9 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M274.21 418.89 L229.99 424.11 L231.32 452.54 L263.72 465.47 L280.83 439.21 L274.21 418.89 Z"
      /><path d="M274.21 418.89 L229.99 424.11 L231.32 452.54 L263.72 465.47 L280.83 439.21 L274.21 418.89 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1091.98 373.07 L1103.05 405.39 L1062.67 422.67 L1040.53 386.28 L1064.61 366.4 L1091.98 373.07 Z"
      /><path d="M1091.98 373.07 L1103.05 405.39 L1062.67 422.67 L1040.53 386.28 L1064.61 366.4 L1091.98 373.07 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M934.54 910.42 L943.35 943.88 L910.29 949.36 L904.8 924.39 L925.65 907.48 L934.54 910.42 Z"
      /><path d="M934.54 910.42 L943.35 943.88 L910.29 949.36 L904.8 924.39 L925.65 907.48 L934.54 910.42 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1513.28 854.83 L1486.12 842.94 L1457.87 871.73 L1478.34 909.48 L1499.6899 907.95 L1521.4399 872.12 L1513.28 854.83 Z"
      /><path d="M1513.28 854.83 L1486.12 842.94 L1457.87 871.73 L1478.34 909.48 L1499.6899 907.95 L1521.4399 872.12 L1513.28 854.83 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1277.4301 594.26 L1276.86 561.7 L1237.75 565.78 L1247.91 605.29 L1277.4301 594.26 Z"
      /><path d="M1277.4301 594.26 L1276.86 561.7 L1237.75 565.78 L1247.91 605.29 L1277.4301 594.26 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M157.58 900.48 L136.4 896.44 L108.59 922.12 L108.34 942.55 L168.96 949.4 L175.39 935 L157.58 900.48 Z"
      /><path d="M157.58 900.48 L136.4 896.44 L108.59 922.12 L108.34 942.55 L168.96 949.4 L175.39 935 L157.58 900.48 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M891.65 326.99 L865.75 361.73 L873.69 377.34 L916.58 381.47 L922.18 340.34 L891.65 326.99 Z"
      /><path d="M891.65 326.99 L865.75 361.73 L873.69 377.34 L916.58 381.47 L922.18 340.34 L891.65 326.99 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1489.09 667.11 L1516.39 697.18 L1513.97 707.88 L1477.71 727.07 L1474.9 726.32 L1457.15 695.82 L1489.09 667.11 Z"
      /><path d="M1489.09 667.11 L1516.39 697.18 L1513.97 707.88 L1477.71 727.07 L1474.9 726.32 L1457.15 695.82 L1489.09 667.11 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M807.29 963.98 L800.46 963.87 L776.45 995.01 L778.2 1016.46 L820.08 1029.89 L852.39 1009.18 L851.48 1006.7 L807.29 963.98 Z"
      /><path d="M807.29 963.98 L800.46 963.87 L776.45 995.01 L778.2 1016.46 L820.08 1029.89 L852.39 1009.18 L851.48 1006.7 L807.29 963.98 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1864.6 370.36 L1897.1801 404.77 L1866.89 439.35 L1857.52 440.85 L1835.27 398.19 L1864.6 370.36 Z"
      /><path d="M1864.6 370.36 L1897.1801 404.77 L1866.89 439.35 L1857.52 440.85 L1835.27 398.19 L1864.6 370.36 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M840.07 679.27 L813.9 707.14 L816.53 728.79 L832.32 740.36 L848.07 737.57 L872.62 702.37 L859.29 680.55 L840.07 679.27 Z"
      /><path d="M840.07 679.27 L813.9 707.14 L816.53 728.79 L832.32 740.36 L848.07 737.57 L872.62 702.37 L859.29 680.55 L840.07 679.27 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M518.77 974.99 L538.09 984.73 L548.42 1006.69 L544.19 1022.5 L507.63 1037.78 L482.74 1017.07 L483.66 994.61 L518.77 974.99 Z"
      /><path d="M518.77 974.99 L538.09 984.73 L548.42 1006.69 L544.19 1022.5 L507.63 1037.78 L482.74 1017.07 L483.66 994.61 L518.77 974.99 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M587.79 853.63 L557.72 850.34 L551.47 854.31 L544.18 887.72 L561.23 907.15 L597.36 898.92 L603.56 889.34 L587.79 853.63 Z"
      /><path d="M587.79 853.63 L557.72 850.34 L551.47 854.31 L544.18 887.72 L561.23 907.15 L597.36 898.92 L603.56 889.34 L587.79 853.63 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M223.3 270.05 L233.19 286.06 L221.27 336.96 L196.63 340.12 L184.49 333.54 L176.21 292.73 L223.3 270.05 Z"
      /><path d="M223.3 270.05 L233.19 286.06 L221.27 336.96 L196.63 340.12 L184.49 333.54 L176.21 292.73 L223.3 270.05 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1163.72 487.98 L1197.17 517.92 L1181.79 545.07 L1160.59 548.29 L1148.63 538.72 L1149.9 495.53 L1163.72 487.98 Z"
      /><path d="M1163.72 487.98 L1197.17 517.92 L1181.79 545.07 L1160.59 548.29 L1148.63 538.72 L1149.9 495.53 L1163.72 487.98 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M400.96 910.48 L374.42 881.95 L345.01 895.39 L343.1 932.3 L386.65 938.23 L400.96 910.48 Z"
      /><path d="M400.96 910.48 L374.42 881.95 L345.01 895.39 L343.1 932.3 L386.65 938.23 L400.96 910.48 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M105.46 946.86 L55.14 947.88 L46.17 974.8 L55.45 991.36 L91.49 995.71 L107.3 976.57 L105.46 946.86 Z"
      /><path d="M105.46 946.86 L55.14 947.88 L46.17 974.8 L55.45 991.36 L91.49 995.71 L107.3 976.57 L105.46 946.86 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1563.1801 975.38 L1519.88 964.62 L1509.52 973.32 L1522.37 1022.36 L1557.78 1024.0601 L1563.1801 975.38 Z"
      /><path d="M1563.1801 975.38 L1519.88 964.62 L1509.52 973.32 L1522.37 1022.36 L1557.78 1024.0601 L1563.1801 975.38 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M483.85 696.09 L536.49 724.49 L537.58 738.54 L514.52 768.4 L475.22 747.21 L468.08 714.33 L483.85 696.09 Z"
      /><path d="M483.85 696.09 L536.49 724.49 L537.58 738.54 L514.52 768.4 L475.22 747.21 L468.08 714.33 L483.85 696.09 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M983.58 1045.48 L958.73 1028.3101 L924.77 1034.8199 L919.3 1080 L984 1080 L983.58 1045.48 Z"
      /><path d="M983.58 1045.48 L958.73 1028.3101 L924.77 1034.8199 L919.3 1080 L984 1080 L983.58 1045.48 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1018.03 328.21 L1022.96 332.49 L1021.63 383.02 L1019.57 383.9 L974.76 366.47 L972.85 354.65 L989.9 329.61 L1018.03 328.21 Z"
      /><path d="M1018.03 328.21 L1022.96 332.49 L1021.63 383.02 L1019.57 383.9 L974.76 366.47 L972.85 354.65 L989.9 329.61 L1018.03 328.21 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M177.38 644.64 L162.59 613 L135.07 618.35 L124.78 637.59 L133.73 655.33 L149.79 661.02 L177.38 644.64 Z"
      /><path d="M177.38 644.64 L162.59 613 L135.07 618.35 L124.78 637.59 L133.73 655.33 L149.79 661.02 L177.38 644.64 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M177.38 644.64 L184.66 647.07 L198.87 684.07 L169.6 703.49 L168.41 703.39 L155.57 693.74 L149.79 661.02 L177.38 644.64 Z"
      /><path d="M177.38 644.64 L184.66 647.07 L198.87 684.07 L169.6 703.49 L168.41 703.39 L155.57 693.74 L149.79 661.02 L177.38 644.64 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1102.59 774.56 L1082.52 750.54 L1042.42 763.01 L1038.34 772.18 L1043.62 789.99 L1074.79 807.8 L1102.59 774.56 Z"
      /><path d="M1102.59 774.56 L1082.52 750.54 L1042.42 763.01 L1038.34 772.18 L1043.62 789.99 L1074.79 807.8 L1102.59 774.56 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1165.23 987.42 L1142.79 946.05 L1121.61 956.78 L1114.84 990.79 L1120.85 998.52 L1135.29 1002.51 L1165.23 987.42 Z"
      /><path d="M1165.23 987.42 L1142.79 946.05 L1121.61 956.78 L1114.84 990.79 L1120.85 998.52 L1135.29 1002.51 L1165.23 987.42 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1495.34 187.86 L1484.6 186.25 L1450.51 231.38 L1483.9399 250.83 L1501.17 245.07 L1513.15 221 L1495.34 187.86 Z"
      /><path d="M1495.34 187.86 L1484.6 186.25 L1450.51 231.38 L1483.9399 250.83 L1501.17 245.07 L1513.15 221 L1495.34 187.86 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1106.39 855.76 L1139.66 868.84 L1141.45 871.64 L1125.88 906.06 L1096.52 907.91 L1086.1 874.92 L1106.39 855.76 Z"
      /><path d="M1106.39 855.76 L1139.66 868.84 L1141.45 871.64 L1125.88 906.06 L1096.52 907.91 L1086.1 874.92 L1106.39 855.76 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1243.64 783.21 L1216.03 763.56 L1192.04 783.43 L1201.51 807.14 L1241.62 798.67 L1243.64 783.21 Z"
      /><path d="M1243.64 783.21 L1216.03 763.56 L1192.04 783.43 L1201.51 807.14 L1241.62 798.67 L1243.64 783.21 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1543.28 503.15 L1521.04 501.48 L1501.65 522.45 L1501.33 538.35 L1520.63 557.13 L1534.17 558.1 L1560.25 538.15 L1562.9399 523.64 L1543.28 503.15 Z"
      /><path d="M1543.28 503.15 L1521.04 501.48 L1501.65 522.45 L1501.33 538.35 L1520.63 557.13 L1534.17 558.1 L1560.25 538.15 L1562.9399 523.64 L1543.28 503.15 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M61.05 505.76 L39.72 514.88 L51.32 547.29 L61.35 546.95 L78.83 519.98 L77.76 515.25 L61.05 505.76 Z"
      /><path d="M61.05 505.76 L39.72 514.88 L51.32 547.29 L61.35 546.95 L78.83 519.98 L77.76 515.25 L61.05 505.76 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M577.13 72.25 L599.39 87.83 L594.41 126.09 L551.01 110.14 L550.41 85.84 L577.13 72.25 Z"
      /><path d="M577.13 72.25 L599.39 87.83 L594.41 126.09 L551.01 110.14 L550.41 85.84 L577.13 72.25 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M988.39 954.11 L1007.98 964.05 L1010.54 988.64 L1001.39 996.75 L966.98 991.76 L960.66 981.97 L988.39 954.11 Z"
      /><path d="M988.39 954.11 L1007.98 964.05 L1010.54 988.64 L1001.39 996.75 L966.98 991.76 L960.66 981.97 L988.39 954.11 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1450.5601 777.54 L1437.89 795.58 L1438.87 810.08 L1482.1 828.76 L1498.96 797.5 L1490.79 779.05 L1450.5601 777.54 Z"
      /><path d="M1450.5601 777.54 L1437.89 795.58 L1438.87 810.08 L1482.1 828.76 L1498.96 797.5 L1490.79 779.05 L1450.5601 777.54 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M280.93 1029.77 L227.84 1014.05 L205.89 1035.39 L204.91 1039.0601 L213.7 1080 L278 1080 L280.93 1029.77 Z"
      /><path d="M280.93 1029.77 L227.84 1014.05 L205.89 1035.39 L204.91 1039.0601 L213.7 1080 L278 1080 L280.93 1029.77 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M55.45 991.36 L91.49 995.71 L99.7 1027.76 L84.25 1044.98 L45.42 1033.74 L40.81 1025.8199 L55.45 991.36 Z"
      /><path d="M55.45 991.36 L91.49 995.71 L99.7 1027.76 L84.25 1044.98 L45.42 1033.74 L40.81 1025.8199 L55.45 991.36 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M602.07 282.65 L570.81 285.57 L564.49 308.4 L592.27 324.09 L611.94 313.77 L614.26 305.08 L602.07 282.65 Z"
      /><path d="M602.07 282.65 L570.81 285.57 L564.49 308.4 L592.27 324.09 L611.94 313.77 L614.26 305.08 L602.07 282.65 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M664.9 0 L665.33 33.02 L678.81 46.7 L720.83 33.46 L721.9 0 L664.9 0 Z"
      /><path d="M664.9 0 L665.33 33.02 L678.81 46.7 L720.83 33.46 L721.9 0 L664.9 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M63.2 625.96 L49.47 619.61 L43.3 622.13 L28.16 653.1 L42.26 668.98 L74.11 664.15 L63.2 625.96 Z"
      /><path d="M63.2 625.96 L49.47 619.61 L43.3 622.13 L28.16 653.1 L42.26 668.98 L74.11 664.15 L63.2 625.96 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M460.19 811.18 L488.41 851.34 L487 855.96 L442.61 882.65 L415.5 841.26 L455.38 809.48 L460.19 811.18 Z"
      /><path d="M460.19 811.18 L488.41 851.34 L487 855.96 L442.61 882.65 L415.5 841.26 L455.38 809.48 L460.19 811.18 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1257.58 339.88 L1240.74 339.55 L1220.09 372.22 L1225.61 386.41 L1250.6899 392.88 L1270.79 364.93 L1257.58 339.88 Z"
      /><path d="M1257.58 339.88 L1240.74 339.55 L1220.09 372.22 L1225.61 386.41 L1250.6899 392.88 L1270.79 364.93 L1257.58 339.88 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1106.86 291.26 L1140.3101 328.1 L1128.03 344.74 L1111.92 347.33 L1088.38 325.73 L1097.03 295.61 L1106.86 291.26 Z"
      /><path d="M1106.86 291.26 L1140.3101 328.1 L1128.03 344.74 L1111.92 347.33 L1088.38 325.73 L1097.03 295.61 L1106.86 291.26 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M938.81 598.18 L949.89 634.62 L921.71 662.31 L892.96 645.49 L905.57 599.27 L938.81 598.18 Z"
      /><path d="M938.81 598.18 L949.89 634.62 L921.71 662.31 L892.96 645.49 L905.57 599.27 L938.81 598.18 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1848.23 292.33 L1825.05 279.94 L1797.85 290.99 L1790.3101 331.65 L1806.29 344.29 L1837.28 337.23 L1848.23 292.33 Z"
      /><path d="M1848.23 292.33 L1825.05 279.94 L1797.85 290.99 L1790.3101 331.65 L1806.29 344.29 L1837.28 337.23 L1848.23 292.33 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M114.41 504.9 L112.73 529.84 L96.83 534.46 L78.83 519.98 L77.76 515.25 L97.23 497.89 L114.41 504.9 Z"
      /><path d="M114.41 504.9 L112.73 529.84 L96.83 534.46 L78.83 519.98 L77.76 515.25 L97.23 497.89 L114.41 504.9 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M605.81 1036.52 L601.86 1034.64 L565.52 1046.7 L560.8 1080 L613.4 1080 L605.81 1036.52 Z"
      /><path d="M605.81 1036.52 L601.86 1034.64 L565.52 1046.7 L560.8 1080 L613.4 1080 L605.81 1036.52 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1417.35 737.13 L1445.17 750.44 L1450.5601 777.54 L1437.89 795.58 L1391.86 774.86 L1391.6 774.3 L1398.35 750.09 L1417.35 737.13 Z"
      /><path d="M1417.35 737.13 L1445.17 750.44 L1450.5601 777.54 L1437.89 795.58 L1391.86 774.86 L1391.6 774.3 L1398.35 750.09 L1417.35 737.13 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1791.05 181.08 L1791.11 181.08 L1806.24 225.52 L1761.73 252.06 L1749.1801 244.76 L1734.53 209.06 L1734.89 208.17 L1791.05 181.08 Z"
      /><path d="M1791.05 181.08 L1791.11 181.08 L1806.24 225.52 L1761.73 252.06 L1749.1801 244.76 L1734.53 209.06 L1734.89 208.17 L1791.05 181.08 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M955.41 186.63 L999.01 194.34 L1003.76 199.86 L998.56 227.28 L967.55 245.97 L952.17 241.84 L932.66 202.83 L955.41 186.63 Z"
      /><path d="M955.41 186.63 L999.01 194.34 L1003.76 199.86 L998.56 227.28 L967.55 245.97 L952.17 241.84 L932.66 202.83 L955.41 186.63 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M228.9 100.96 L238.02 106.29 L231.25 157.86 L228.02 160.6 L200.66 156.85 L181.95 120.71 L187.92 111.21 L228.9 100.96 Z"
      /><path d="M228.9 100.96 L238.02 106.29 L231.25 157.86 L228.02 160.6 L200.66 156.85 L181.95 120.71 L187.92 111.21 L228.9 100.96 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M780.64 887.05 L739.65 893.02 L730.06 908.77 L742.53 939.37 L781.72 937.38 L792.56 901.89 L780.64 887.05 Z"
      /><path d="M780.64 887.05 L739.65 893.02 L730.06 908.77 L742.53 939.37 L781.72 937.38 L792.56 901.89 L780.64 887.05 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1911.01 157.27 L1920 158.2 L1920 226.4 L1875.01 228.34 L1861.79 218.72 L1860.7 183.37 L1911.01 157.27 Z"
      /><path d="M1911.01 157.27 L1920 158.2 L1920 226.4 L1875.01 228.34 L1861.79 218.72 L1860.7 183.37 L1911.01 157.27 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1523.41 320.71 L1521.74 319.76 L1482.8 338.56 L1480.24 362.57 L1515.95 374.92 L1530.04 358.66 L1523.41 320.71 Z"
      /><path d="M1523.41 320.71 L1521.74 319.76 L1482.8 338.56 L1480.24 362.57 L1515.95 374.92 L1530.04 358.66 L1523.41 320.71 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1255.01 820.63 L1256.99 821.28 L1274.61 849.34 L1268.97 868.47 L1227.04 871.53 L1225.79 870.02 L1225.73 842.92 L1255.01 820.63 Z"
      /><path d="M1255.01 820.63 L1256.99 821.28 L1274.61 849.34 L1268.97 868.47 L1227.04 871.53 L1225.79 870.02 L1225.73 842.92 L1255.01 820.63 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1066.9399 244.95 L1065.58 283.38 L1056.35 290.69 L1023.43 288.52 L1016.47 280.2 L1022.73 251.74 L1063.83 239.39 L1066.9399 244.95 Z"
      /><path d="M1066.9399 244.95 L1065.58 283.38 L1056.35 290.69 L1023.43 288.52 L1016.47 280.2 L1022.73 251.74 L1063.83 239.39 L1066.9399 244.95 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M141.94 817.71 L119.69 804.35 L99.61 809.61 L90.25 850.42 L95.87 858.52 L122.35 863.2 L145.99 841.22 L141.94 817.71 Z"
      /><path d="M141.94 817.71 L119.69 804.35 L99.61 809.61 L90.25 850.42 L95.87 858.52 L122.35 863.2 L145.99 841.22 L141.94 817.71 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M143.49 572.87 L129.31 572.72 L118.5 594.74 L135.07 618.35 L162.59 613 L168.17 600.87 L143.49 572.87 Z"
      /><path d="M143.49 572.87 L129.31 572.72 L118.5 594.74 L135.07 618.35 L162.59 613 L168.17 600.87 L143.49 572.87 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1225.61 386.41 L1250.6899 392.88 L1262.85 415.31 L1249.37 437.67 L1220.26 440.25 L1201.66 415.02 L1225.61 386.41 Z"
      /><path d="M1225.61 386.41 L1250.6899 392.88 L1262.85 415.31 L1249.37 437.67 L1220.26 440.25 L1201.66 415.02 L1225.61 386.41 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M441.66 412.86 L422.51 386.7 L395.18 387.43 L386.27 398.57 L388.43 423.74 L418.39 439.75 L430.58 434.5 L441.66 412.86 Z"
      /><path d="M441.66 412.86 L422.51 386.7 L395.18 387.43 L386.27 398.57 L388.43 423.74 L418.39 439.75 L430.58 434.5 L441.66 412.86 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1592.5 568.56 L1569.71 597.76 L1555.04 597.2 L1534.17 558.1 L1560.25 538.15 L1592.5 568.56 Z"
      /><path d="M1592.5 568.56 L1569.71 597.76 L1555.04 597.2 L1534.17 558.1 L1560.25 538.15 L1592.5 568.56 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M571.75 636.2 L546.15 642.13 L536.57 668.57 L556.45 692.3 L585.45 662.54 L576.14 638.19 L571.75 636.2 Z"
      /><path d="M571.75 636.2 L546.15 642.13 L536.57 668.57 L556.45 692.3 L585.45 662.54 L576.14 638.19 L571.75 636.2 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M921.12 989.13 L920.4 1029.73 L866.53 1022.19 L856.7 1011.05 L905.6 976.68 L921.12 989.13 Z"
      /><path d="M921.12 989.13 L920.4 1029.73 L866.53 1022.19 L856.7 1011.05 L905.6 976.68 L921.12 989.13 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1143.8 810.8 L1136.13 809.13 L1102.12 833.08 L1106.39 855.76 L1139.66 868.84 L1152.78 822.52 L1143.8 810.8 Z"
      /><path d="M1143.8 810.8 L1136.13 809.13 L1102.12 833.08 L1106.39 855.76 L1139.66 868.84 L1152.78 822.52 L1143.8 810.8 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1143.95 206.5 L1175.3199 222.58 L1176.76 241.35 L1138.6801 265.9 L1124.89 262.55 L1123.7 221.51 L1143.95 206.5 Z"
      /><path d="M1143.95 206.5 L1175.3199 222.58 L1176.76 241.35 L1138.6801 265.9 L1124.89 262.55 L1123.7 221.51 L1143.95 206.5 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1264.63 465.53 L1249.37 437.67 L1220.26 440.25 L1209.3199 465.89 L1223.7 488.04 L1254.5 484.83 L1264.63 465.53 Z"
      /><path d="M1264.63 465.53 L1249.37 437.67 L1220.26 440.25 L1209.3199 465.89 L1223.7 488.04 L1254.5 484.83 L1264.63 465.53 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1857.67 1020.59 L1877.12 1039.75 L1874.4 1080 L1826.1 1080 L1824.39 1044.76 L1852.9 1020.41 L1857.67 1020.59 Z"
      /><path d="M1857.67 1020.59 L1877.12 1039.75 L1874.4 1080 L1826.1 1080 L1824.39 1044.76 L1852.9 1020.41 L1857.67 1020.59 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M198.4 0 L204.34 47.76 L221.2 55.86 L256.9 41.73 L258.1 0 L198.4 0 Z"
      /><path d="M198.4 0 L204.34 47.76 L221.2 55.86 L256.9 41.73 L258.1 0 L198.4 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1378.96 569.67 L1342.1801 559.61 L1320.98 582.33 L1320.11 591.87 L1344.36 612.57 L1361.48 608.27 L1378.96 569.67 Z"
      /><path d="M1378.96 569.67 L1342.1801 559.61 L1320.98 582.33 L1320.11 591.87 L1344.36 612.57 L1361.48 608.27 L1378.96 569.67 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1712.4 0 L1771.3 0 L1773.5601 18.05 L1750.5 54.93 L1735.46 55.24 L1711.63 36.59 L1712.4 0 Z"
      /><path d="M1712.4 0 L1771.3 0 L1773.5601 18.05 L1750.5 54.93 L1735.46 55.24 L1711.63 36.59 L1712.4 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M592.27 324.09 L588.98 351.69 L564.58 365.39 L554.79 359.3 L555.82 313.01 L564.49 308.4 L592.27 324.09 Z"
      /><path d="M592.27 324.09 L588.98 351.69 L564.58 365.39 L554.79 359.3 L555.82 313.01 L564.49 308.4 L592.27 324.09 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1090.9399 208.97 L1123.7 221.51 L1124.89 262.55 L1122.62 263.84 L1066.9399 244.95 L1063.83 239.39 L1065.25 231.04 L1090.9399 208.97 Z"
      /><path d="M1090.9399 208.97 L1123.7 221.51 L1124.89 262.55 L1122.62 263.84 L1066.9399 244.95 L1063.83 239.39 L1065.25 231.04 L1090.9399 208.97 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M98.49 168.81 L138.53 182.88 L126.47 231.31 L111.83 234.5 L80.89 211.7 L88.28 176.88 L98.49 168.81 Z"
      /><path d="M98.49 168.81 L138.53 182.88 L126.47 231.31 L111.83 234.5 L80.89 211.7 L88.28 176.88 L98.49 168.81 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M609.89 33.14 L578.64 45.89 L577.13 72.25 L599.39 87.83 L626.47 76.3 L626.81 47.71 L609.89 33.14 Z"
      /><path d="M609.89 33.14 L578.64 45.89 L577.13 72.25 L599.39 87.83 L626.47 76.3 L626.81 47.71 L609.89 33.14 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M92.84 267.22 L54.22 261.12 L45.17 274.73 L47.72 304.12 L84.46 313.33 L104.94 298.43 L92.84 267.22 Z"
      /><path d="M92.84 267.22 L54.22 261.12 L45.17 274.73 L47.72 304.12 L84.46 313.33 L104.94 298.43 L92.84 267.22 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M118.5 594.74 L135.07 618.35 L124.78 637.59 L104.42 636.37 L89.96 617.71 L95.85 599.58 L118.5 594.74 Z"
      /><path d="M118.5 594.74 L135.07 618.35 L124.78 637.59 L104.42 636.37 L89.96 617.71 L95.85 599.58 L118.5 594.74 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1324.33 307.61 L1308.17 327.93 L1313.59 351.51 L1346.84 357.43 L1364.64 335.87 L1359.61 316.26 L1324.33 307.61 Z"
      /><path d="M1324.33 307.61 L1308.17 327.93 L1313.59 351.51 L1346.84 357.43 L1364.64 335.87 L1359.61 316.26 L1324.33 307.61 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1341.9 71.49 L1331.58 107.63 L1303.9301 110.89 L1285.26 93.47 L1283.64 85.19 L1319 56.45 L1341.9 71.49 Z"
      /><path d="M1341.9 71.49 L1331.58 107.63 L1303.9301 110.89 L1285.26 93.47 L1283.64 85.19 L1319 56.45 L1341.9 71.49 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1426 826.41 L1380.27 823.74 L1379.0601 824.62 L1375.4399 852.93 L1386.0699 868.1 L1426.4399 872.21 L1431.71 868.3 L1426 826.41 Z"
      /><path d="M1426 826.41 L1380.27 823.74 L1379.0601 824.62 L1375.4399 852.93 L1386.0699 868.1 L1426.4399 872.21 L1431.71 868.3 L1426 826.41 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M28.16 653.1 L42.26 668.98 L34.75 699.43 L0 698.2 L0 654.4 L28.16 653.1 Z"
      /><path d="M28.16 653.1 L42.26 668.98 L34.75 699.43 L0 698.2 L0 654.4 L28.16 653.1 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1739.13 835.86 L1752.73 843.92 L1756.09 895.2 L1741.7 907.94 L1718.8 904.56 L1699.75 868.54 L1739.13 835.86 Z"
      /><path d="M1739.13 835.86 L1752.73 843.92 L1756.09 895.2 L1741.7 907.94 L1718.8 904.56 L1699.75 868.54 L1739.13 835.86 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1397.6 89.62 L1382.48 91.62 L1362.1899 123.16 L1380.61 142.51 L1406.36 137.63 L1405.9399 98.43 L1397.6 89.62 Z"
      /><path d="M1397.6 89.62 L1382.48 91.62 L1362.1899 123.16 L1380.61 142.51 L1406.36 137.63 L1405.9399 98.43 L1397.6 89.62 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M274.35 79.86 L239.96 106.08 L277.99 130.71 L301.14 106.97 L301.85 103.1 L274.35 79.86 Z"
      /><path d="M274.35 79.86 L239.96 106.08 L277.99 130.71 L301.14 106.97 L301.85 103.1 L274.35 79.86 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M635.26 337.81 L623.43 366.86 L588.98 351.69 L592.27 324.09 L611.94 313.77 L635.26 337.81 Z"
      /><path d="M635.26 337.81 L623.43 366.86 L588.98 351.69 L592.27 324.09 L611.94 313.77 L635.26 337.81 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M469.37 317.29 L487.76 345.7 L465.77 368.46 L439.12 360.82 L431.35 340.3 L468.69 317.27 L469.37 317.29 Z"
      /><path d="M469.37 317.29 L487.76 345.7 L465.77 368.46 L439.12 360.82 L431.35 340.3 L468.69 317.27 L469.37 317.29 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1453.72 440.9 L1473.84 476.71 L1463.17 496.76 L1459.6801 498.15 L1427.52 482.81 L1425.3101 457.51 L1444.3101 437.91 L1453.72 440.9 Z"
      /><path d="M1453.72 440.9 L1473.84 476.71 L1463.17 496.76 L1459.6801 498.15 L1427.52 482.81 L1425.3101 457.51 L1444.3101 437.91 L1453.72 440.9 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M884.6 849.77 L922.93 857.6 L925.76 866.67 L916.75 886.74 L879.52 890.79 L879.04 890.19 L884.6 849.77 Z"
      /><path d="M884.6 849.77 L922.93 857.6 L925.76 866.67 L916.75 886.74 L879.52 890.79 L879.04 890.19 L884.6 849.77 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M440.49 488.16 L409.91 473.91 L396.73 480.86 L393.26 515.78 L433.22 528.29 L440.27 520.9 L440.49 488.16 Z"
      /><path d="M440.49 488.16 L409.91 473.91 L396.73 480.86 L393.26 515.78 L433.22 528.29 L440.27 520.9 L440.49 488.16 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M0 1020.1 L40.81 1025.8199 L45.42 1033.74 L30.3 1080 L0 1080 L0 1020.1 Z"
      /><path d="M0 1020.1 L40.81 1025.8199 L45.42 1033.74 L30.3 1080 L0 1080 L0 1020.1 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1790.8 447.52 L1757.6 447.79 L1734.78 491.62 L1760.46 508.52 L1791.53 503.05 L1802.42 459.56 L1790.8 447.52 Z"
      /><path d="M1790.8 447.52 L1757.6 447.79 L1734.78 491.62 L1760.46 508.52 L1791.53 503.05 L1802.42 459.56 L1790.8 447.52 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1043.62 789.99 L1018.94 822.52 L988.57 809.73 L993.28 773.63 L1038.34 772.18 L1043.62 789.99 Z"
      /><path d="M1043.62 789.99 L1018.94 822.52 L988.57 809.73 L993.28 773.63 L1038.34 772.18 L1043.62 789.99 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1566.46 826.17 L1567.92 866.89 L1552.27 879.72 L1521.4399 872.12 L1513.28 854.83 L1545.12 818.14 L1566.46 826.17 Z"
      /><path d="M1566.46 826.17 L1567.92 866.89 L1552.27 879.72 L1521.4399 872.12 L1513.28 854.83 L1545.12 818.14 L1566.46 826.17 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M757.95 703.32 L739.87 699.1 L726.63 704.85 L716.54 737.73 L735.26 763.18 L770.76 756.84 L775.8 745.34 L757.95 703.32 Z"
      /><path d="M757.95 703.32 L739.87 699.1 L726.63 704.85 L716.54 737.73 L735.26 763.18 L770.76 756.84 L775.8 745.34 L757.95 703.32 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1102.12 833.08 L1077.47 818.44 L1051.78 847.65 L1060.09 869.56 L1086.1 874.92 L1106.39 855.76 L1102.12 833.08 Z"
      /><path d="M1102.12 833.08 L1077.47 818.44 L1051.78 847.65 L1060.09 869.56 L1086.1 874.92 L1106.39 855.76 L1102.12 833.08 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1286.88 22.57 L1316.4 44.46 L1319 56.45 L1283.64 85.19 L1259.03 66.54 L1256.41 55.33 L1286.88 22.57 Z"
      /><path d="M1286.88 22.57 L1316.4 44.46 L1319 56.45 L1283.64 85.19 L1259.03 66.54 L1256.41 55.33 L1286.88 22.57 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M770.4 33.42 L790.42 45.49 L793.01 61.65 L766.51 84.35 L736.7 55.72 L736.55 50.62 L770.4 33.42 Z"
      /><path d="M770.4 33.42 L790.42 45.49 L793.01 61.65 L766.51 84.35 L736.7 55.72 L736.55 50.62 L770.4 33.42 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M693.22 855.86 L726.59 858.11 L739.65 893.02 L730.06 908.77 L698.88 908.65 L684.8 881.69 L693.22 855.86 Z"
      /><path d="M693.22 855.86 L726.59 858.11 L739.65 893.02 L730.06 908.77 L698.88 908.65 L684.8 881.69 L693.22 855.86 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1579.85 423.74 L1596.2 432.19 L1596.64 433.25 L1586.1 472.56 L1559.33 468.3 L1547.35 451.51 L1579.85 423.74 Z"
      /><path d="M1579.85 423.74 L1596.2 432.19 L1596.64 433.25 L1586.1 472.56 L1559.33 468.3 L1547.35 451.51 L1579.85 423.74 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1026.5699 50.18 L1010.44 94.13 L1022.56 109.96 L1058.45 102.17 L1070.41 63.91 L1066.78 58.68 L1026.5699 50.18 Z"
      /><path d="M1026.5699 50.18 L1010.44 94.13 L1022.56 109.96 L1058.45 102.17 L1070.41 63.91 L1066.78 58.68 L1026.5699 50.18 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M312.83 591.24 L312.53 608.53 L280.97 629.96 L267.22 620.04 L262.99 589.74 L290.11 574.14 L312.83 591.24 Z"
      /><path d="M312.83 591.24 L312.53 608.53 L280.97 629.96 L267.22 620.04 L262.99 589.74 L290.11 574.14 L312.83 591.24 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M892.96 645.49 L921.71 662.31 L927.54 688.37 L892.13 707.66 L872.62 702.37 L859.29 680.55 L877.51 649.41 L892.96 645.49 Z"
      /><path d="M892.96 645.49 L921.71 662.31 L927.54 688.37 L892.13 707.66 L872.62 702.37 L859.29 680.55 L877.51 649.41 L892.96 645.49 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1447.5601 592.15 L1418.15 562.85 L1392.65 570.82 L1413.87 623.79 L1423.52 626.58 L1447.5601 592.15 Z"
      /><path d="M1447.5601 592.15 L1418.15 562.85 L1392.65 570.82 L1413.87 623.79 L1423.52 626.58 L1447.5601 592.15 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M723.43 543.07 L710.88 571.75 L695.36 575.01 L671.28 558.67 L670.14 550.3 L706.84 524.28 L723.43 543.07 Z"
      /><path d="M723.43 543.07 L710.88 571.75 L695.36 575.01 L671.28 558.67 L670.14 550.3 L706.84 524.28 L723.43 543.07 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M56.19 900.29 L44 926.65 L0 927 L0 874 L34.29 872.34 L56.19 900.29 Z"
      /><path d="M56.19 900.29 L44 926.65 L0 927 L0 874 L34.29 872.34 L56.19 900.29 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1423.52 626.58 L1413.87 623.79 L1386.5699 630.94 L1370.24 666.27 L1372.29 677.95 L1379.4301 685.07 L1428.92 662.82 L1433.1 642.15 L1423.52 626.58 Z"
      /><path d="M1423.52 626.58 L1413.87 623.79 L1386.5699 630.94 L1370.24 666.27 L1372.29 677.95 L1379.4301 685.07 L1428.92 662.82 L1433.1 642.15 L1423.52 626.58 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1798.15 120.87 L1753.01 118.95 L1752.36 119.35 L1748.7 144.97 L1791.05 181.08 L1791.11 181.08 L1802.0699 170.98 L1798.15 120.87 Z"
      /><path d="M1798.15 120.87 L1753.01 118.95 L1752.36 119.35 L1748.7 144.97 L1791.05 181.08 L1791.11 181.08 L1802.0699 170.98 L1798.15 120.87 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1261.79 639.1 L1252.58 634.16 L1223.02 660.41 L1246.33 684.2 L1272.05 674.12 L1261.79 639.1 Z"
      /><path d="M1261.79 639.1 L1252.58 634.16 L1223.02 660.41 L1246.33 684.2 L1272.05 674.12 L1261.79 639.1 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M560.5 523.59 L565.74 546.27 L528.58 567.54 L522.54 560.83 L522.64 523.84 L541.1 512.38 L560.5 523.59 Z"
      /><path d="M560.5 523.59 L565.74 546.27 L528.58 567.54 L522.54 560.83 L522.64 523.84 L541.1 512.38 L560.5 523.59 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M40.4 117 L0 115.4 L0 163.6 L41.19 166.46 L42.56 165.33 L49.25 130.53 L40.4 117 Z"
      /><path d="M40.4 117 L0 115.4 L0 163.6 L41.19 166.46 L42.56 165.33 L49.25 130.53 L40.4 117 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M972.75 524.19 L1000.48 552.85 L984.45 585.74 L947.93 587.73 L939.23 541.11 L972.75 524.19 Z"
      /><path d="M972.75 524.19 L1000.48 552.85 L984.45 585.74 L947.93 587.73 L939.23 541.11 L972.75 524.19 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M655.9 294.31 L656.1 330.73 L635.26 337.81 L611.94 313.77 L614.26 305.08 L650.55 288.65 L655.9 294.31 Z"
      /><path d="M655.9 294.31 L656.1 330.73 L635.26 337.81 L611.94 313.77 L614.26 305.08 L650.55 288.65 L655.9 294.31 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1026.5699 50.18 L1019.25 40.41 L981.49 43.76 L966.81 77.92 L975.02 89.76 L1010.44 94.13 L1026.5699 50.18 Z"
      /><path d="M1026.5699 50.18 L1019.25 40.41 L981.49 43.76 L966.81 77.92 L975.02 89.76 L1010.44 94.13 L1026.5699 50.18 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1586.36 768.71 L1547.01 774.53 L1536.91 803.11 L1545.12 818.14 L1566.46 826.17 L1575.05 822.53 L1595.08 781.59 L1586.36 768.71 Z"
      /><path d="M1586.36 768.71 L1547.01 774.53 L1536.91 803.11 L1545.12 818.14 L1566.46 826.17 L1575.05 822.53 L1595.08 781.59 L1586.36 768.71 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M764.33 575.07 L746.84 543.03 L723.43 543.07 L710.88 571.75 L736.25 598.88 L737.16 599.01 L764.33 575.07 Z"
      /><path d="M764.33 575.07 L746.84 543.03 L723.43 543.07 L710.88 571.75 L736.25 598.88 L737.16 599.01 L764.33 575.07 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M880.93 828.16 L881.74 845.78 L835.41 859.21 L821.69 842.89 L841.43 814.2 L880.93 828.16 Z"
      /><path d="M880.93 828.16 L881.74 845.78 L835.41 859.21 L821.69 842.89 L841.43 814.2 L880.93 828.16 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M205.17 530.29 L207.19 534.83 L200.98 553.18 L183.88 559.66 L164.51 551.15 L156.76 525.29 L166.66 515.86 L175.66 513.11 L205.17 530.29 Z"
      /><path d="M205.17 530.29 L207.19 534.83 L200.98 553.18 L183.88 559.66 L164.51 551.15 L156.76 525.29 L166.66 515.86 L175.66 513.11 L205.17 530.29 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M439.9 212.21 L442.9 226.34 L402.77 250.57 L388.62 243.38 L385.96 213.95 L402.33 197.04 L439.9 212.21 Z"
      /><path d="M439.9 212.21 L442.9 226.34 L402.77 250.57 L388.62 243.38 L385.96 213.95 L402.33 197.04 L439.9 212.21 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1571.35 700.37 L1540.0699 684.66 L1516.39 697.18 L1513.97 707.88 L1535.12 737.48 L1567.24 723.3 L1571.35 700.37 Z"
      /><path d="M1571.35 700.37 L1540.0699 684.66 L1516.39 697.18 L1513.97 707.88 L1535.12 737.48 L1567.24 723.3 L1571.35 700.37 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1855.74 766.8 L1827.27 761.98 L1799.89 789.56 L1804.5601 812.33 L1846.54 830.24 L1857.02 826.37 L1867.73 802.62 L1855.74 766.8 Z"
      /><path d="M1855.74 766.8 L1827.27 761.98 L1799.89 789.56 L1804.5601 812.33 L1846.54 830.24 L1857.02 826.37 L1867.73 802.62 L1855.74 766.8 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M716.65 997.86 L720.88 1024.34 L690.73 1036.8 L670.31 1013.63 L670.24 1004.04 L683.13 990.41 L716.65 997.86 Z"
      /><path d="M716.65 997.86 L720.88 1024.34 L690.73 1036.8 L670.31 1013.63 L670.24 1004.04 L683.13 990.41 L716.65 997.86 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M267.39 337.98 L271.25 342.21 L263.92 382.07 L236.45 382.13 L225.26 339.52 L267.39 337.98 Z"
      /><path d="M267.39 337.98 L271.25 342.21 L263.92 382.07 L236.45 382.13 L225.26 339.52 L267.39 337.98 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1920 403.4 L1920 473.8 L1866.89 439.35 L1897.1801 404.77 L1920 403.4 Z"
      /><path d="M1920 403.4 L1920 473.8 L1866.89 439.35 L1897.1801 404.77 L1920 403.4 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1675.8 394.9 L1649.03 433.26 L1620.51 405.76 L1620.84 386.35 L1675.8 394.9 Z"
      /><path d="M1675.8 394.9 L1649.03 433.26 L1620.51 405.76 L1620.84 386.35 L1675.8 394.9 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1198.21 591.18 L1163.71 598.67 L1160.4 631.16 L1197.45 643.4 L1212.8101 612.6 L1198.21 591.18 Z"
      /><path d="M1198.21 591.18 L1163.71 598.67 L1160.4 631.16 L1197.45 643.4 L1212.8101 612.6 L1198.21 591.18 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M205.89 1035.39 L156.71 995.54 L154.41 996.65 L135.54 1032.78 L145.1 1053.28 L204.91 1039.0601 L205.89 1035.39 Z"
      /><path d="M205.89 1035.39 L156.71 995.54 L154.41 996.65 L135.54 1032.78 L145.1 1053.28 L204.91 1039.0601 L205.89 1035.39 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1694.4301 217.74 L1671.1899 194.81 L1643.22 201.78 L1644.85 246.27 L1682.8101 257.5 L1694.4301 217.74 Z"
      /><path d="M1694.4301 217.74 L1671.1899 194.81 L1643.22 201.78 L1644.85 246.27 L1682.8101 257.5 L1694.4301 217.74 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M835.03 518.61 L849.66 546.38 L838.49 573.12 L795.53 574.95 L798.01 524.54 L835.03 518.61 Z"
      /><path d="M835.03 518.61 L849.66 546.38 L838.49 573.12 L795.53 574.95 L798.01 524.54 L835.03 518.61 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1920 158.2 L1920 85.1 L1875.45 105.09 L1870.74 118.59 L1911.01 157.27 L1920 158.2 Z"
      /><path d="M1920 158.2 L1920 85.1 L1875.45 105.09 L1870.74 118.59 L1911.01 157.27 L1920 158.2 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M465.97 579.83 L498.36 605.97 L501.58 621.08 L497 628.24 L456.22 640.31 L442.38 605.9 L465.97 579.83 Z"
      /><path d="M465.97 579.83 L498.36 605.97 L501.58 621.08 L497 628.24 L456.22 640.31 L442.38 605.9 L465.97 579.83 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M732.54 412.78 L758.64 418.47 L760.99 451.67 L728.78 472.97 L709.51 457.91 L709.1 432.51 L732.54 412.78 Z"
      /><path d="M732.54 412.78 L758.64 418.47 L760.99 451.67 L728.78 472.97 L709.51 457.91 L709.1 432.51 L732.54 412.78 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M709.51 457.91 L728.78 472.97 L730.05 487.62 L705.64 514.71 L678.31 499.37 L671.49 474.05 L673.34 470.67 L709.51 457.91 Z"
      /><path d="M709.51 457.91 L728.78 472.97 L730.05 487.62 L705.64 514.71 L678.31 499.37 L671.49 474.05 L673.34 470.67 L709.51 457.91 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1021.63 383.02 L1040.53 386.28 L1062.67 422.67 L1054.6 446.76 L1001.96 440.1 L996.72 430.99 L1019.57 383.9 L1021.63 383.02 Z"
      /><path d="M1021.63 383.02 L1040.53 386.28 L1062.67 422.67 L1054.6 446.76 L1001.96 440.1 L996.72 430.99 L1019.57 383.9 L1021.63 383.02 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M542.12 260.95 L526.08 273.91 L522.95 305.37 L524.92 308.38 L555.82 313.01 L564.49 308.4 L570.81 285.57 L562.23 269.05 L542.12 260.95 Z"
      /><path d="M542.12 260.95 L526.08 273.91 L522.95 305.37 L524.92 308.38 L555.82 313.01 L564.49 308.4 L570.81 285.57 L562.23 269.05 L542.12 260.95 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1883.42 848.34 L1857.02 826.37 L1846.54 830.24 L1830.8 872.28 L1862.74 897.73 L1877.5699 887.77 L1883.42 848.34 Z"
      /><path d="M1883.42 848.34 L1857.02 826.37 L1846.54 830.24 L1830.8 872.28 L1862.74 897.73 L1877.5699 887.77 L1883.42 848.34 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1373.36 37.18 L1397.16 43.26 L1407 62.76 L1397.6 89.62 L1382.48 91.62 L1351.62 69.64 L1373.36 37.18 Z"
      /><path d="M1373.36 37.18 L1397.16 43.26 L1407 62.76 L1397.6 89.62 L1382.48 91.62 L1351.62 69.64 L1373.36 37.18 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M807.17 841.91 L784.79 801.16 L745.77 819.34 L745.6 836.99 L783.91 860.82 L807.17 841.91 Z"
      /><path d="M807.17 841.91 L784.79 801.16 L745.77 819.34 L745.6 836.99 L783.91 860.82 L807.17 841.91 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1709.9301 766.03 L1689.51 804.28 L1680.6 807.24 L1646.51 772.51 L1648.48 763.49 L1695.37 741.63 L1709.9301 766.03 Z"
      /><path d="M1709.9301 766.03 L1689.51 804.28 L1680.6 807.24 L1646.51 772.51 L1648.48 763.49 L1695.37 741.63 L1709.9301 766.03 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1920 565 L1920 638.8 L1875.21 637.64 L1870.65 633.44 L1863.85 580.03 L1873.28 568.3 L1920 565 Z"
      /><path d="M1920 565 L1920 638.8 L1875.21 637.64 L1870.65 633.44 L1863.85 580.03 L1873.28 568.3 L1920 565 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M410.23 114.44 L380.48 116.2 L376.64 135.05 L396.22 168.86 L400.17 170.57 L416.78 159.49 L410.23 114.44 Z"
      /><path d="M410.23 114.44 L380.48 116.2 L376.64 135.05 L396.22 168.86 L400.17 170.57 L416.78 159.49 L410.23 114.44 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1783.37 949.91 L1752.3199 943.73 L1733.3101 965.82 L1737.09 990.94 L1789.36 995.88 L1792.27 992.16 L1783.37 949.91 Z"
      /><path d="M1783.37 949.91 L1752.3199 943.73 L1733.3101 965.82 L1737.09 990.94 L1789.36 995.88 L1792.27 992.16 L1783.37 949.91 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1283.78 895.05 L1293.51 912.83 L1277.67 948.72 L1249.76 941.95 L1239.89 915.02 L1283.78 895.05 Z"
      /><path d="M1283.78 895.05 L1293.51 912.83 L1277.67 948.72 L1249.76 941.95 L1239.89 915.02 L1283.78 895.05 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1346.24 123.13 L1331.92 154.05 L1353.24 175.79 L1368.79 174.57 L1380.61 142.51 L1362.1899 123.16 L1346.24 123.13 Z"
      /><path d="M1346.24 123.13 L1331.92 154.05 L1353.24 175.79 L1368.79 174.57 L1380.61 142.51 L1362.1899 123.16 L1346.24 123.13 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M934.04 334.2 L972.85 354.65 L974.76 366.47 L959.35 386.96 L918.25 383.69 L916.58 381.47 L922.18 340.34 L934.04 334.2 Z"
      /><path d="M934.04 334.2 L972.85 354.65 L974.76 366.47 L959.35 386.96 L918.25 383.69 L916.58 381.47 L922.18 340.34 L934.04 334.2 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M414.86 281.7 L383.11 302.43 L406.71 337.52 L424.82 336.66 L425.82 285.88 L414.86 281.7 Z"
      /><path d="M414.86 281.7 L383.11 302.43 L406.71 337.52 L424.82 336.66 L425.82 285.88 L414.86 281.7 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1042.42 763.01 L1028.98 725.99 L989.82 726.69 L982.78 734.49 L983.45 762.21 L993.28 773.63 L1038.34 772.18 L1042.42 763.01 Z"
      /><path d="M1042.42 763.01 L1028.98 725.99 L989.82 726.69 L982.78 734.49 L983.45 762.21 L993.28 773.63 L1038.34 772.18 L1042.42 763.01 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M396.73 480.86 L366.76 467.25 L345.91 484.61 L354.28 521.07 L379.05 526.24 L393.26 515.78 L396.73 480.86 Z"
      /><path d="M396.73 480.86 L366.76 467.25 L345.91 484.61 L354.28 521.07 L379.05 526.24 L393.26 515.78 L396.73 480.86 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M198.87 684.07 L169.6 703.49 L192.91 741.55 L216.28 745.45 L225.8 733.01 L210.79 687.05 L198.87 684.07 Z"
      /><path d="M198.87 684.07 L169.6 703.49 L192.91 741.55 L216.28 745.45 L225.8 733.01 L210.79 687.05 L198.87 684.07 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M527.64 70.85 L502.88 86.18 L504.47 119.59 L530.38 131.69 L551.01 110.14 L550.41 85.84 L527.64 70.85 Z"
      /><path d="M527.64 70.85 L502.88 86.18 L504.47 119.59 L530.38 131.69 L551.01 110.14 L550.41 85.84 L527.64 70.85 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M245.73 207.9 L248.71 245.48 L223.36 269.56 L189.18 226.2 L191.62 216.34 L233.12 200.09 L245.73 207.9 Z"
      /><path d="M245.73 207.9 L248.71 245.48 L223.36 269.56 L189.18 226.2 L191.62 216.34 L233.12 200.09 L245.73 207.9 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1212.8101 612.6 L1197.45 643.4 L1204.87 659.79 L1223.02 660.41 L1252.58 634.16 L1243.72 613.08 L1212.8101 612.6 Z"
      /><path d="M1212.8101 612.6 L1197.45 643.4 L1204.87 659.79 L1223.02 660.41 L1252.58 634.16 L1243.72 613.08 L1212.8101 612.6 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M599.07 602.77 L602.99 622.43 L576.14 638.19 L571.75 636.2 L563.53 596.4 L575.39 590.19 L599.07 602.77 Z"
      /><path d="M599.07 602.77 L602.99 622.43 L576.14 638.19 L571.75 636.2 L563.53 596.4 L575.39 590.19 L599.07 602.77 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M685.56 125.49 L647.77 120.49 L643.93 158.54 L653.69 168.06 L680.37 164.51 L686.77 127.14 L685.56 125.49 Z"
      /><path d="M685.56 125.49 L647.77 120.49 L643.93 158.54 L653.69 168.06 L680.37 164.51 L686.77 127.14 L685.56 125.49 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M322.74 801.23 L342.21 821.47 L341.86 836.34 L318.17 858.37 L283.98 847.14 L281.04 842.75 L287.2 816.13 L322.74 801.23 Z"
      /><path d="M322.74 801.23 L342.21 821.47 L341.86 836.34 L318.17 858.37 L283.98 847.14 L281.04 842.75 L287.2 816.13 L322.74 801.23 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1382.34 447.77 L1376.49 451.74 L1396.39 505.84 L1396.9399 505.85 L1427.52 482.81 L1425.3101 457.51 L1382.34 447.77 Z"
      /><path d="M1382.34 447.77 L1376.49 451.74 L1396.39 505.84 L1396.9399 505.85 L1427.52 482.81 L1425.3101 457.51 L1382.34 447.77 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1103.05 405.39 L1117.8199 411.87 L1126.67 433.27 L1105.99 468.44 L1061.63 461.44 L1054.6 446.76 L1062.67 422.67 L1103.05 405.39 Z"
      /><path d="M1103.05 405.39 L1117.8199 411.87 L1126.67 433.27 L1105.99 468.44 L1061.63 461.44 L1054.6 446.76 L1062.67 422.67 L1103.05 405.39 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M147.24 178.46 L174.56 185.23 L191.62 216.34 L189.18 226.2 L151.41 246.97 L126.47 231.31 L138.53 182.88 L147.24 178.46 Z"
      /><path d="M147.24 178.46 L174.56 185.23 L191.62 216.34 L189.18 226.2 L151.41 246.97 L126.47 231.31 L138.53 182.88 L147.24 178.46 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1509.52 973.32 L1486.05 973.14 L1464.26 992.39 L1461.7 1021.32 L1505.8101 1037.59 L1522.37 1022.36 L1509.52 973.32 Z"
      /><path d="M1509.52 973.32 L1486.05 973.14 L1464.26 992.39 L1461.7 1021.32 L1505.8101 1037.59 L1522.37 1022.36 L1509.52 973.32 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1920 347.8 L1887.2 345.36 L1865.73 359.89 L1864.6 370.36 L1897.1801 404.77 L1920 403.4 L1920 347.8 Z"
      /><path d="M1920 347.8 L1887.2 345.36 L1865.73 359.89 L1864.6 370.36 L1897.1801 404.77 L1920 403.4 L1920 347.8 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M781.72 937.38 L800.46 963.87 L776.45 995.01 L733.75 973.92 L731.17 960.2 L742.53 939.37 L781.72 937.38 Z"
      /><path d="M781.72 937.38 L800.46 963.87 L776.45 995.01 L733.75 973.92 L731.17 960.2 L742.53 939.37 L781.72 937.38 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1129.22 162.93 L1143.4 177.01 L1143.95 206.5 L1123.7 221.51 L1090.9399 208.97 L1089.84 179.95 L1129.22 162.93 Z"
      /><path d="M1129.22 162.93 L1143.4 177.01 L1143.95 206.5 L1123.7 221.51 L1090.9399 208.97 L1089.84 179.95 L1129.22 162.93 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1599.76 874.16 L1609 888.68 L1605.0699 907.6 L1570.7 923.06 L1559.99 917.44 L1552.27 879.72 L1567.92 866.89 L1599.76 874.16 Z"
      /><path d="M1599.76 874.16 L1609 888.68 L1605.0699 907.6 L1570.7 923.06 L1559.99 917.44 L1552.27 879.72 L1567.92 866.89 L1599.76 874.16 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1024.46 838.68 L1051.78 847.65 L1060.09 869.56 L1041.4 893.66 L1019.48 885.18 L1005.97 862.02 L1024.46 838.68 Z"
      /><path d="M1024.46 838.68 L1051.78 847.65 L1060.09 869.56 L1041.4 893.66 L1019.48 885.18 L1005.97 862.02 L1024.46 838.68 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M360.15 35.1 L379.28 61.24 L371 73.63 L328.15 78.14 L316.26 44.51 L360.15 35.1 Z"
      /><path d="M360.15 35.1 L379.28 61.24 L371 73.63 L328.15 78.14 L316.26 44.51 L360.15 35.1 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M570.89 952.7 L556.12 931.42 L515.88 941.16 L518.77 974.99 L538.09 984.73 L570.89 952.7 Z"
      /><path d="M570.89 952.7 L556.12 931.42 L515.88 941.16 L518.77 974.99 L538.09 984.73 L570.89 952.7 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M733.23 356.72 L768.9 367.18 L769.89 409.54 L758.64 418.47 L732.54 412.78 L720 385.76 L733.23 356.72 Z"
      /><path d="M733.23 356.72 L768.9 367.18 L769.89 409.54 L758.64 418.47 L732.54 412.78 L720 385.76 L733.23 356.72 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1205.77 570.4 L1181.79 545.07 L1160.59 548.29 L1152.26 586.65 L1163.71 598.67 L1198.21 591.18 L1205.77 570.4 Z"
      /><path d="M1205.77 570.4 L1181.79 545.07 L1160.59 548.29 L1152.26 586.65 L1163.71 598.67 L1198.21 591.18 L1205.77 570.4 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M318.17 858.37 L323.48 883.01 L284.66 912.01 L279.61 911.81 L269.44 896.61 L283.98 847.14 L318.17 858.37 Z"
      /><path d="M318.17 858.37 L323.48 883.01 L284.66 912.01 L279.61 911.81 L269.44 896.61 L283.98 847.14 L318.17 858.37 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1216.34 748 L1198.74 729.21 L1189.37 729.57 L1166.59 764.65 L1171 775.25 L1192.04 783.43 L1216.03 763.56 L1216.34 748 Z"
      /><path d="M1216.34 748 L1198.74 729.21 L1189.37 729.57 L1166.59 764.65 L1171 775.25 L1192.04 783.43 L1216.03 763.56 L1216.34 748 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1754.4301 557.35 L1801.72 558.53 L1814.04 583.98 L1801.49 611.6 L1746.54 602.05 L1741.4 567.52 L1754.4301 557.35 Z"
      /><path d="M1754.4301 557.35 L1801.72 558.53 L1814.04 583.98 L1801.49 611.6 L1746.54 602.05 L1741.4 567.52 L1754.4301 557.35 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1061.63 461.44 L1105.99 468.44 L1115.64 488.17 L1093.9399 527.93 L1089.5 528.79 L1044.89 502.75 L1061.63 461.44 Z"
      /><path d="M1061.63 461.44 L1105.99 468.44 L1115.64 488.17 L1093.9399 527.93 L1089.5 528.79 L1044.89 502.75 L1061.63 461.44 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M893.09 546.65 L894.65 590.01 L852.86 597.26 L838.49 573.12 L849.66 546.38 L893.09 546.65 Z"
      /><path d="M893.09 546.65 L894.65 590.01 L852.86 597.26 L838.49 573.12 L849.66 546.38 L893.09 546.65 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M628.58 1029.45 L605.81 1036.52 L613.4 1080 L644.6 1080 L652.1 1054.14 L643.02 1035.6899 L628.58 1029.45 Z"
      /><path d="M628.58 1029.45 L605.81 1036.52 L613.4 1080 L644.6 1080 L652.1 1054.14 L643.02 1035.6899 L628.58 1029.45 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1418.35 145.5 L1406.36 137.63 L1380.61 142.51 L1368.79 174.57 L1384.04 187.96 L1426.0699 175.24 L1426.51 174.53 L1418.35 145.5 Z"
      /><path d="M1418.35 145.5 L1406.36 137.63 L1380.61 142.51 L1368.79 174.57 L1384.04 187.96 L1426.0699 175.24 L1426.51 174.53 L1418.35 145.5 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1682.91 1039.1801 L1674.46 1015.79 L1640.92 1016.11 L1634.17 1041.53 L1665.23 1063.58 L1682.91 1039.1801 Z"
      /><path d="M1682.91 1039.1801 L1674.46 1015.79 L1640.92 1016.11 L1634.17 1041.53 L1665.23 1063.58 L1682.91 1039.1801 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M200.66 156.85 L174.56 185.23 L147.24 178.46 L150.18 128.19 L181.95 120.71 L200.66 156.85 Z"
      /><path d="M200.66 156.85 L174.56 185.23 L147.24 178.46 L150.18 128.19 L181.95 120.71 L200.66 156.85 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M903.14 44.85 L884.22 69.05 L855.28 66.81 L845.28 54.12 L844.4 41.76 L848.55 34.88 L892.55 25.16 L903.14 44.85 Z"
      /><path d="M903.14 44.85 L884.22 69.05 L855.28 66.81 L845.28 54.12 L844.4 41.76 L848.55 34.88 L892.55 25.16 L903.14 44.85 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M684.67 826.87 L647.05 797.98 L622.13 828.84 L641.24 851.76 L684.07 842.62 L684.67 826.87 Z"
      /><path d="M684.67 826.87 L647.05 797.98 L622.13 828.84 L641.24 851.76 L684.07 842.62 L684.67 826.87 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M745.46 222.01 L771.31 225.5 L776.4 231.33 L771.09 263.35 L749.06 275.39 L731.42 250.36 L736.44 228.16 L745.46 222.01 Z"
      /><path d="M745.46 222.01 L771.31 225.5 L776.4 231.33 L771.09 263.35 L749.06 275.39 L731.42 250.36 L736.44 228.16 L745.46 222.01 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1627.83 727.63 L1648.48 763.49 L1646.51 772.51 L1621.48 788.64 L1595.08 781.59 L1586.36 768.71 L1589.4399 748.92 L1627.83 727.63 Z"
      /><path d="M1627.83 727.63 L1648.48 763.49 L1646.51 772.51 L1621.48 788.64 L1595.08 781.59 L1586.36 768.71 L1589.4399 748.92 L1627.83 727.63 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M693.69 175.91 L702.6 176.55 L715.04 191.51 L709.84 216.41 L699.68 221.61 L674.46 211.8 L693.69 175.91 Z"
      /><path d="M693.69 175.91 L702.6 176.55 L715.04 191.51 L709.84 216.41 L699.68 221.61 L674.46 211.8 L693.69 175.91 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1533.52 431.66 L1543.2 449.96 L1509.12 471.17 L1501.39 467.72 L1493.74 425.22 L1494.96 423.23 L1533.52 431.66 Z"
      /><path d="M1533.52 431.66 L1543.2 449.96 L1509.12 471.17 L1501.39 467.72 L1493.74 425.22 L1494.96 423.23 L1533.52 431.66 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M553.65 436.87 L532.67 447.06 L523.72 474.55 L541 489.5 L574.44 474.38 L553.65 436.87 Z"
      /><path d="M553.65 436.87 L532.67 447.06 L523.72 474.55 L541 489.5 L574.44 474.38 L553.65 436.87 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1682.01 565.16 L1674.3199 592.24 L1639.47 607.83 L1632.8199 605.32 L1610.71 565.86 L1622.1801 548.17 L1644.62 544.08 L1682.01 565.16 Z"
      /><path d="M1682.01 565.16 L1674.3199 592.24 L1639.47 607.83 L1632.8199 605.32 L1610.71 565.86 L1622.1801 548.17 L1644.62 544.08 L1682.01 565.16 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1694.4 951.34 L1733.3101 965.82 L1737.09 990.94 L1728.53 1004.45 L1684.95 998.44 L1677.02 971.5 L1694.4 951.34 Z"
      /><path d="M1694.4 951.34 L1733.3101 965.82 L1737.09 990.94 L1728.53 1004.45 L1684.95 998.44 L1677.02 971.5 L1694.4 951.34 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M320.99 324.12 L354.79 348.54 L340.74 376.24 L308.51 369.58 L301 346.71 L320.99 324.12 Z"
      /><path d="M320.99 324.12 L354.79 348.54 L340.74 376.24 L308.51 369.58 L301 346.71 L320.99 324.12 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1615.59 699.49 L1576.27 697.03 L1571.35 700.37 L1567.24 723.3 L1589.4399 748.92 L1627.83 727.63 L1630.04 717.57 L1615.59 699.49 Z"
      /><path d="M1615.59 699.49 L1576.27 697.03 L1571.35 700.37 L1567.24 723.3 L1589.4399 748.92 L1627.83 727.63 L1630.04 717.57 L1615.59 699.49 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1306.09 395.11 L1340.59 403.63 L1343.2 443.54 L1307.8199 451.9 L1288.99 415.46 L1306.09 395.11 Z"
      /><path d="M1306.09 395.11 L1340.59 403.63 L1343.2 443.54 L1307.8199 451.9 L1288.99 415.46 L1306.09 395.11 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1609.1801 379.36 L1617.1801 380.46 L1620.84 386.35 L1620.51 405.76 L1596.2 432.19 L1579.85 423.74 L1571.2 403.82 L1609.1801 379.36 Z"
      /><path d="M1609.1801 379.36 L1617.1801 380.46 L1620.84 386.35 L1620.51 405.76 L1596.2 432.19 L1579.85 423.74 L1571.2 403.82 L1609.1801 379.36 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1501.65 522.45 L1463.17 496.76 L1459.6801 498.15 L1443.35 534.39 L1470.66 552.84 L1501.33 538.35 L1501.65 522.45 Z"
      /><path d="M1501.65 522.45 L1463.17 496.76 L1459.6801 498.15 L1443.35 534.39 L1470.66 552.84 L1501.33 538.35 L1501.65 522.45 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M121.15 728.44 L144.66 735.18 L156.91 761.78 L125.76 773.69 L105.54 755.78 L115.21 730.98 L121.15 728.44 Z"
      /><path d="M121.15 728.44 L144.66 735.18 L156.91 761.78 L125.76 773.69 L105.54 755.78 L115.21 730.98 L121.15 728.44 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1615.3101 837.22 L1575.05 822.53 L1566.46 826.17 L1567.92 866.89 L1599.76 874.16 L1615.3101 837.22 Z"
      /><path d="M1615.3101 837.22 L1575.05 822.53 L1566.46 826.17 L1567.92 866.89 L1599.76 874.16 L1615.3101 837.22 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1501.39 467.72 L1473.84 476.71 L1453.72 440.9 L1493.74 425.22 L1501.39 467.72 Z"
      /><path d="M1501.39 467.72 L1473.84 476.71 L1453.72 440.9 L1493.74 425.22 L1501.39 467.72 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M783.91 860.82 L745.6 836.99 L726.59 858.11 L739.65 893.02 L780.64 887.05 L783.91 860.82 Z"
      /><path d="M783.91 860.82 L745.6 836.99 L726.59 858.11 L739.65 893.02 L780.64 887.05 L783.91 860.82 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M545.98 407.82 L513.66 398.05 L503.77 428.49 L532.67 447.06 L553.65 436.87 L553.73 436.71 L545.98 407.82 Z"
      /><path d="M545.98 407.82 L513.66 398.05 L503.77 428.49 L532.67 447.06 L553.65 436.87 L553.73 436.71 L545.98 407.82 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1137.3199 62.67 L1129.74 61.72 L1112.25 72.32 L1108.73 120.16 L1128.9399 134.34 L1160.98 117.95 L1165.5699 97.6 L1137.3199 62.67 Z"
      /><path d="M1137.3199 62.67 L1129.74 61.72 L1112.25 72.32 L1108.73 120.16 L1128.9399 134.34 L1160.98 117.95 L1165.5699 97.6 L1137.3199 62.67 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M468.69 317.27 L431.35 340.3 L424.82 336.66 L425.82 285.88 L433.6 284.63 L468.69 317.27 Z"
      /><path d="M468.69 317.27 L431.35 340.3 L424.82 336.66 L425.82 285.88 L433.6 284.63 L468.69 317.27 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M229.99 424.11 L231.32 452.54 L217.26 464.71 L175.38 445.92 L175.47 444.2 L216.17 408.5 L229.99 424.11 Z"
      /><path d="M229.99 424.11 L231.32 452.54 L217.26 464.71 L175.38 445.92 L175.47 444.2 L216.17 408.5 L229.99 424.11 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M574.27 221.62 L587.74 234.41 L587.95 243.66 L562.23 269.05 L542.12 260.95 L540.2 247.17 L555.64 222.82 L574.27 221.62 Z"
      /><path d="M574.27 221.62 L587.74 234.41 L587.95 243.66 L562.23 269.05 L542.12 260.95 L540.2 247.17 L555.64 222.82 L574.27 221.62 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1033.46 678.97 L1040.3101 709.93 L1028.98 725.99 L989.82 726.69 L984.42 680.39 L986.05 677.94 L1033.46 678.97 Z"
      /><path d="M1033.46 678.97 L1040.3101 709.93 L1028.98 725.99 L989.82 726.69 L984.42 680.39 L986.05 677.94 L1033.46 678.97 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M345.01 895.39 L323.48 883.01 L284.66 912.01 L328.45 945.09 L343.1 932.3 L345.01 895.39 Z"
      /><path d="M345.01 895.39 L323.48 883.01 L284.66 912.01 L328.45 945.09 L343.1 932.3 L345.01 895.39 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1432.09 0.23 L1455.37 59.71 L1455.34 59.75 L1407 62.76 L1397.16 43.26 L1432.09 0.23 Z"
      /><path d="M1432.09 0.23 L1455.37 59.71 L1455.34 59.75 L1407 62.76 L1397.16 43.26 L1432.09 0.23 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M407.8 0 L403.41 58.07 L415.43 64.45 L445.52 55.89 L440.8 0 L407.8 0 Z"
      /><path d="M407.8 0 L403.41 58.07 L415.43 64.45 L445.52 55.89 L440.8 0 L407.8 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M535.58 198.25 L502.95 224.37 L540.2 247.17 L555.64 222.82 L535.58 198.25 Z"
      /><path d="M535.58 198.25 L502.95 224.37 L540.2 247.17 L555.64 222.82 L535.58 198.25 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M694.49 657.67 L661.1 653.16 L651.03 673 L656.87 700.93 L664.09 707.68 L698.45 689.56 L694.49 657.67 Z"
      /><path d="M694.49 657.67 L661.1 653.16 L651.03 673 L656.87 700.93 L664.09 707.68 L698.45 689.56 L694.49 657.67 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1737.1899 830.44 L1689.51 804.28 L1680.6 807.24 L1670.9301 823.76 L1689.72 866.49 L1699.75 868.54 L1739.13 835.86 L1737.1899 830.44 Z"
      /><path d="M1737.1899 830.44 L1689.51 804.28 L1680.6 807.24 L1670.9301 823.76 L1689.72 866.49 L1699.75 868.54 L1739.13 835.86 L1737.1899 830.44 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M551.47 854.31 L513.68 839.55 L488.41 851.34 L487 855.96 L508.77 895.99 L544.18 887.72 L551.47 854.31 Z"
      /><path d="M551.47 854.31 L513.68 839.55 L488.41 851.34 L487 855.96 L508.77 895.99 L544.18 887.72 L551.47 854.31 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M85.3 433.9 L84.67 467.94 L61.76 476.13 L42.96 467.45 L39.1 438.29 L74.18 426.98 L85.3 433.9 Z"
      /><path d="M85.3 433.9 L84.67 467.94 L61.76 476.13 L42.96 467.45 L39.1 438.29 L74.18 426.98 L85.3 433.9 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M665.14 738.08 L670.4 745.89 L668.55 764 L646.99 788.19 L593.81 762.4 L593.53 760.72 L604.66 738.71 L665.14 738.08 Z"
      /><path d="M665.14 738.08 L670.4 745.89 L668.55 764 L646.99 788.19 L593.81 762.4 L593.53 760.72 L604.66 738.71 L665.14 738.08 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1461.7 1021.32 L1505.8101 1037.59 L1507 1080 L1450.9 1080 L1447.71 1032.67 L1461.7 1021.32 Z"
      /><path d="M1461.7 1021.32 L1505.8101 1037.59 L1507 1080 L1450.9 1080 L1447.71 1032.67 L1461.7 1021.32 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M617.88 629.23 L621.76 640.02 L610.54 669.6 L610.52 669.61 L585.45 662.54 L576.14 638.19 L602.99 622.43 L617.88 629.23 Z"
      /><path d="M617.88 629.23 L621.76 640.02 L610.54 669.6 L610.52 669.61 L585.45 662.54 L576.14 638.19 L602.99 622.43 L617.88 629.23 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M872.62 702.37 L848.07 737.57 L883.46 764.73 L903.34 752.27 L892.13 707.66 L872.62 702.37 Z"
      /><path d="M872.62 702.37 L848.07 737.57 L883.46 764.73 L903.34 752.27 L892.13 707.66 L872.62 702.37 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1339.49 224.66 L1378.5601 229.68 L1381.8199 277.55 L1325.02 265.41 L1339.49 224.66 Z"
      /><path d="M1339.49 224.66 L1378.5601 229.68 L1381.8199 277.55 L1325.02 265.41 L1339.49 224.66 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M474 0 L440.8 0 L445.52 55.89 L466.45 64 L486.19 37.92 L474 0 Z"
      /><path d="M474 0 L440.8 0 L445.52 55.89 L466.45 64 L486.19 37.92 L474 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M61.76 476.13 L42.96 467.45 L20.62 483.83 L35.48 513.66 L39.72 514.88 L61.05 505.76 L61.76 476.13 Z"
      /><path d="M61.76 476.13 L42.96 467.45 L20.62 483.83 L35.48 513.66 L39.72 514.88 L61.05 505.76 L61.76 476.13 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M440.55 713.32 L413.76 752.58 L417.28 767.92 L441.63 778.47 L475.22 747.21 L468.08 714.33 L440.55 713.32 Z"
      /><path d="M440.55 713.32 L413.76 752.58 L417.28 767.92 L441.63 778.47 L475.22 747.21 L468.08 714.33 L440.55 713.32 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M95.87 858.52 L122.35 863.2 L136.4 896.44 L108.59 922.12 L78.39 895.87 L95.87 858.52 Z"
      /><path d="M95.87 858.52 L122.35 863.2 L136.4 896.44 L108.59 922.12 L78.39 895.87 L95.87 858.52 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1718.8 904.56 L1691.83 929.7 L1694.4 951.34 L1733.3101 965.82 L1752.3199 943.73 L1741.7 907.94 L1718.8 904.56 Z"
      /><path d="M1718.8 904.56 L1691.83 929.7 L1694.4 951.34 L1733.3101 965.82 L1752.3199 943.73 L1741.7 907.94 L1718.8 904.56 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1734.53 209.06 L1749.1801 244.76 L1705.15 270.66 L1686.13 263.57 L1682.8101 257.5 L1694.4301 217.74 L1734.53 209.06 Z"
      /><path d="M1734.53 209.06 L1749.1801 244.76 L1705.15 270.66 L1686.13 263.57 L1682.8101 257.5 L1694.4301 217.74 L1734.53 209.06 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M408.31 840.08 L377.79 862.57 L341.86 836.34 L342.21 821.47 L384.54 799.66 L408.31 840.08 Z"
      /><path d="M408.31 840.08 L377.79 862.57 L341.86 836.34 L342.21 821.47 L384.54 799.66 L408.31 840.08 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M224.75 984.05 L227.84 1014.05 L205.89 1035.39 L156.71 995.54 L172.22 969.16 L224.75 984.05 Z"
      /><path d="M224.75 984.05 L227.84 1014.05 L205.89 1035.39 L156.71 995.54 L172.22 969.16 L224.75 984.05 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1520.63 557.13 L1534.17 558.1 L1555.04 597.2 L1532.5699 616.7 L1498.28 598.89 L1520.63 557.13 Z"
      /><path d="M1520.63 557.13 L1534.17 558.1 L1555.04 597.2 L1532.5699 616.7 L1498.28 598.89 L1520.63 557.13 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M176.21 292.73 L184.49 333.54 L143.75 349.94 L136.95 347.25 L121.68 302.89 L155.2 281.85 L176.21 292.73 Z"
      /><path d="M176.21 292.73 L184.49 333.54 L143.75 349.94 L136.95 347.25 L121.68 302.89 L155.2 281.85 L176.21 292.73 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1521.4399 872.12 L1552.27 879.72 L1559.99 917.44 L1524.03 932.1 L1499.6899 907.95 L1521.4399 872.12 Z"
      /><path d="M1521.4399 872.12 L1552.27 879.72 L1559.99 917.44 L1524.03 932.1 L1499.6899 907.95 L1521.4399 872.12 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1852.28 518.53 L1873.28 568.3 L1863.85 580.03 L1814.04 583.98 L1801.72 558.53 L1813.6801 525.98 L1852.28 518.53 Z"
      /><path d="M1852.28 518.53 L1873.28 568.3 L1863.85 580.03 L1814.04 583.98 L1801.72 558.53 L1813.6801 525.98 L1852.28 518.53 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M808.7 0 L844.9 0 L848.55 34.88 L844.4 41.76 L808.99 29.99 L808.7 0 Z"
      /><path d="M808.7 0 L844.9 0 L848.55 34.88 L844.4 41.76 L808.99 29.99 L808.7 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1089.38 673.18 L1044.83 662.1 L1033.46 678.97 L1040.3101 709.93 L1080.78 714.46 L1089.38 673.18 Z"
      /><path d="M1089.38 673.18 L1044.83 662.1 L1033.46 678.97 L1040.3101 709.93 L1080.78 714.46 L1089.38 673.18 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M474 0 L522.1 0 L517.93 37.77 L486.19 37.92 L474 0 Z"
      /><path d="M474 0 L522.1 0 L517.93 37.77 L486.19 37.92 L474 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1300.75 462.61 L1264.63 465.53 L1254.5 484.83 L1272.59 517.93 L1308.88 494.76 L1300.75 462.61 Z"
      /><path d="M1300.75 462.61 L1264.63 465.53 L1254.5 484.83 L1272.59 517.93 L1308.88 494.76 L1300.75 462.61 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1842.1899 459.25 L1858.72 507.52 L1852.28 518.53 L1813.6801 525.98 L1791.53 503.05 L1802.42 459.56 L1842.1899 459.25 Z"
      /><path d="M1842.1899 459.25 L1858.72 507.52 L1852.28 518.53 L1813.6801 525.98 L1791.53 503.05 L1802.42 459.56 L1842.1899 459.25 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M789.63 788.62 L770.76 756.84 L735.26 763.18 L720.96 795.79 L745.77 819.34 L784.79 801.16 L789.63 788.62 Z"
      /><path d="M789.63 788.62 L770.76 756.84 L735.26 763.18 L720.96 795.79 L745.77 819.34 L784.79 801.16 L789.63 788.62 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M931.45 690.81 L927.54 688.37 L892.13 707.66 L903.34 752.27 L922.52 755.08 L944.61 727.04 L931.45 690.81 Z"
      /><path d="M931.45 690.81 L927.54 688.37 L892.13 707.66 L903.34 752.27 L922.52 755.08 L944.61 727.04 L931.45 690.81 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M0 163.6 L0 202.7 L30.86 206.87 L38.77 201.36 L41.19 166.46 L0 163.6 Z"
      /><path d="M0 163.6 L0 202.7 L30.86 206.87 L38.77 201.36 L41.19 166.46 L0 163.6 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1455.34 59.75 L1448.14 100.48 L1405.9399 98.43 L1397.6 89.62 L1407 62.76 L1455.34 59.75 Z"
      /><path d="M1455.34 59.75 L1448.14 100.48 L1405.9399 98.43 L1397.6 89.62 L1407 62.76 L1455.34 59.75 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M536.57 668.57 L508.44 668.63 L483.88 695.82 L483.85 696.09 L536.49 724.49 L556.73 695.47 L556.45 692.3 L536.57 668.57 Z"
      /><path d="M536.57 668.57 L508.44 668.63 L483.88 695.82 L483.85 696.09 L536.49 724.49 L556.73 695.47 L556.45 692.3 L536.57 668.57 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M498.24 224.93 L482.01 181.42 L456.13 184.28 L439.9 212.21 L442.9 226.34 L450.27 232.61 L494.34 229.32 L498.24 224.93 Z"
      /><path d="M498.24 224.93 L482.01 181.42 L456.13 184.28 L439.9 212.21 L442.9 226.34 L450.27 232.61 L494.34 229.32 L498.24 224.93 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1083.6 0 L1066.78 58.68 L1026.5699 50.18 L1019.25 40.41 L1024.6 0 L1083.6 0 Z"
      /><path d="M1083.6 0 L1066.78 58.68 L1026.5699 50.18 L1019.25 40.41 L1024.6 0 L1083.6 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M593.53 760.72 L593.81 762.4 L581.58 791.17 L559.85 801.51 L522.86 790.57 L515.71 781.42 L514.52 768.4 L537.58 738.54 L593.53 760.72 Z"
      /><path d="M593.53 760.72 L593.81 762.4 L581.58 791.17 L559.85 801.51 L522.86 790.57 L515.71 781.42 L514.52 768.4 L537.58 738.54 L593.53 760.72 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M306.74 662.91 L284.04 650.54 L254.45 675.29 L265.77 700.95 L307.49 703.68 L315.31 692.92 L306.74 662.91 Z"
      /><path d="M306.74 662.91 L284.04 650.54 L254.45 675.29 L265.77 700.95 L307.49 703.68 L315.31 692.92 L306.74 662.91 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M583.44 189.71 L566.1 175.01 L536.15 192.35 L535.58 198.25 L555.64 222.82 L574.27 221.62 L583.44 189.71 Z"
      /><path d="M583.44 189.71 L566.1 175.01 L536.15 192.35 L535.58 198.25 L555.64 222.82 L574.27 221.62 L583.44 189.71 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1315.73 838.9 L1294.11 799.68 L1256.99 821.28 L1274.61 849.34 L1315.73 838.9 Z"
      /><path d="M1315.73 838.9 L1294.11 799.68 L1256.99 821.28 L1274.61 849.34 L1315.73 838.9 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M79.98 581.27 L95.85 599.58 L89.96 617.71 L63.2 625.96 L49.47 619.61 L54.32 589.83 L79.98 581.27 Z"
      /><path d="M79.98 581.27 L95.85 599.58 L89.96 617.71 L63.2 625.96 L49.47 619.61 L54.32 589.83 L79.98 581.27 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1328.86 865.23 L1283.85 894.29 L1283.78 895.05 L1293.51 912.83 L1326.5601 922.09 L1343.6899 900.13 L1329.34 865.52 L1328.86 865.23 Z"
      /><path d="M1328.86 865.23 L1283.85 894.29 L1283.78 895.05 L1293.51 912.83 L1326.5601 922.09 L1343.6899 900.13 L1329.34 865.52 L1328.86 865.23 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M647.01 119.64 L647.77 120.49 L643.93 158.54 L614.45 162.96 L594.21 134.31 L595.02 127.31 L647.01 119.64 Z"
      /><path d="M647.01 119.64 L647.77 120.49 L643.93 158.54 L614.45 162.96 L594.21 134.31 L595.02 127.31 L647.01 119.64 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1852.9 1020.41 L1824.39 1044.76 L1788.9399 1026.83 L1789.36 995.88 L1792.27 992.16 L1826.09 986.92 L1852.9 1020.41 Z"
      /><path d="M1852.9 1020.41 L1824.39 1044.76 L1788.9399 1026.83 L1789.36 995.88 L1792.27 992.16 L1826.09 986.92 L1852.9 1020.41 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1338.6 510.38 L1308.88 494.76 L1272.59 517.93 L1272.52 518.23 L1286.72 547.47 L1331.91 531.87 L1338.6 510.38 Z"
      /><path d="M1338.6 510.38 L1308.88 494.76 L1272.59 517.93 L1272.52 518.23 L1286.72 547.47 L1331.91 531.87 L1338.6 510.38 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M901.98 163.58 L886.75 162.05 L864.47 182.76 L864.67 209.5 L894.37 223.33 L928.41 202.01 L901.98 163.58 Z"
      /><path d="M901.98 163.58 L886.75 162.05 L864.47 182.76 L864.67 209.5 L894.37 223.33 L928.41 202.01 L901.98 163.58 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M922.52 755.08 L903.34 752.27 L883.46 764.73 L879.6 777.64 L894.66 809.32 L922.21 809.48 L937.97 792.54 L939.1 779.31 L922.52 755.08 Z"
      /><path d="M922.52 755.08 L903.34 752.27 L883.46 764.73 L879.6 777.64 L894.66 809.32 L922.21 809.48 L937.97 792.54 L939.1 779.31 L922.52 755.08 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M84.25 1044.98 L45.42 1033.74 L30.3 1080 L88.1 1080 L84.25 1044.98 Z"
      /><path d="M84.25 1044.98 L45.42 1033.74 L30.3 1080 L88.1 1080 L84.25 1044.98 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1450.51 231.38 L1483.9399 250.83 L1476.26 287.07 L1455.78 299.92 L1428.72 265.91 L1439.97 232.47 L1450.51 231.38 Z"
      /><path d="M1450.51 231.38 L1483.9399 250.83 L1476.26 287.07 L1455.78 299.92 L1428.72 265.91 L1439.97 232.47 L1450.51 231.38 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M0 744.3 L18.75 746.32 L36.14 777.41 L0 800.1 L0 744.3 Z"
      /><path d="M0 744.3 L18.75 746.32 L36.14 777.41 L0 800.1 L0 744.3 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1237.75 565.78 L1247.91 605.29 L1243.72 613.08 L1212.8101 612.6 L1198.21 591.18 L1205.77 570.4 L1231.6801 561.6 L1237.75 565.78 Z"
      /><path d="M1237.75 565.78 L1247.91 605.29 L1243.72 613.08 L1212.8101 612.6 L1198.21 591.18 L1205.77 570.4 L1231.6801 561.6 L1237.75 565.78 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M570.89 952.7 L573.21 953.46 L590.69 995.21 L590.03 996.39 L548.42 1006.69 L538.09 984.73 L570.89 952.7 Z"
      /><path d="M570.89 952.7 L573.21 953.46 L590.69 995.21 L590.03 996.39 L548.42 1006.69 L538.09 984.73 L570.89 952.7 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M819.05 213.36 L851.83 218.36 L848.98 261.93 L820.75 264.69 L807.56 229.46 L819.05 213.36 Z"
      /><path d="M819.05 213.36 L851.83 218.36 L848.98 261.93 L820.75 264.69 L807.56 229.46 L819.05 213.36 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M158.3 0 L198.4 0 L204.34 47.76 L171.93 65.17 L153.48 60.47 L146.04 44.13 L158.3 0 Z"
      /><path d="M158.3 0 L198.4 0 L204.34 47.76 L171.93 65.17 L153.48 60.47 L146.04 44.13 L158.3 0 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M615.81 984.44 L590.69 995.21 L573.21 953.46 L609.15 941.82 L615.81 984.44 Z"
      /><path d="M615.81 984.44 L590.69 995.21 L573.21 953.46 L609.15 941.82 L615.81 984.44 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1344.36 612.57 L1334.5601 639.57 L1313.95 648.22 L1294.51 627.32 L1296.55 606.25 L1320.11 591.87 L1344.36 612.57 Z"
      /><path d="M1344.36 612.57 L1334.5601 639.57 L1313.95 648.22 L1294.51 627.32 L1296.55 606.25 L1320.11 591.87 L1344.36 612.57 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M37.52 390.99 L68.52 391.71 L74.18 426.98 L39.1 438.29 L26.73 429.83 L37.52 390.99 Z"
      /><path d="M37.52 390.99 L68.52 391.71 L74.18 426.98 L39.1 438.29 L26.73 429.83 L37.52 390.99 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1197.45 643.4 L1160.4 631.16 L1147.47 640.99 L1143.8199 667.87 L1170.48 685.41 L1197.38 673.94 L1204.87 659.79 L1197.45 643.4 Z"
      /><path d="M1197.45 643.4 L1160.4 631.16 L1147.47 640.99 L1143.8199 667.87 L1170.48 685.41 L1197.38 673.94 L1204.87 659.79 L1197.45 643.4 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1704.73 628.04 L1674.3199 592.24 L1639.47 607.83 L1647.38 652.72 L1671.25 664.74 L1677.38 663.45 L1704.73 628.04 Z"
      /><path d="M1704.73 628.04 L1674.3199 592.24 L1639.47 607.83 L1647.38 652.72 L1671.25 664.74 L1677.38 663.45 L1704.73 628.04 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1121.61 956.78 L1092.38 944.08 L1070.26 977.26 L1081.6801 989.5 L1114.84 990.79 L1121.61 956.78 Z"
      /><path d="M1121.61 956.78 L1092.38 944.08 L1070.26 977.26 L1081.6801 989.5 L1114.84 990.79 L1121.61 956.78 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1520.63 557.13 L1501.33 538.35 L1470.66 552.84 L1466.65 588.2 L1486.66 601.61 L1498.28 598.89 L1520.63 557.13 Z"
      /><path d="M1520.63 557.13 L1501.33 538.35 L1470.66 552.84 L1466.65 588.2 L1486.66 601.61 L1498.28 598.89 L1520.63 557.13 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1284.02 773.12 L1258.17 771.4 L1243.64 783.21 L1241.62 798.67 L1255.01 820.63 L1256.99 821.28 L1294.11 799.68 L1297.38 787.42 L1284.02 773.12 Z"
      /><path d="M1284.02 773.12 L1258.17 771.4 L1243.64 783.21 L1241.62 798.67 L1255.01 820.63 L1256.99 821.28 L1294.11 799.68 L1297.38 787.42 L1284.02 773.12 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1860.4301 694.84 L1871.98 704 L1872.36 751.89 L1855.74 766.8 L1827.27 761.98 L1812.29 724.29 L1841.14 696.19 L1860.4301 694.84 Z"
      /><path d="M1860.4301 694.84 L1871.98 704 L1872.36 751.89 L1855.74 766.8 L1827.27 761.98 L1812.29 724.29 L1841.14 696.19 L1860.4301 694.84 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M917.6 274.59 L917.95 274.61 L944.58 302.65 L934.04 334.2 L922.18 340.34 L891.65 326.99 L885.38 311.33 L917.6 274.59 Z"
      /><path d="M917.6 274.59 L917.95 274.61 L944.58 302.65 L934.04 334.2 L922.18 340.34 L891.65 326.99 L885.38 311.33 L917.6 274.59 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1023.43 288.52 L1056.35 290.69 L1058.8101 331.92 L1022.96 332.49 L1018.03 328.21 L1023.43 288.52 Z"
      /><path d="M1023.43 288.52 L1056.35 290.69 L1058.8101 331.92 L1022.96 332.49 L1018.03 328.21 L1023.43 288.52 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1649 879.35 L1609 888.68 L1605.0699 907.6 L1631.9301 936.44 L1661.99 914.45 L1658.83 884.39 L1649 879.35 Z"
      /><path d="M1649 879.35 L1609 888.68 L1605.0699 907.6 L1631.9301 936.44 L1661.99 914.45 L1658.83 884.39 L1649 879.35 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M912.11 485.86 L872.73 446.1 L840.16 473.4 L845.17 497.66 L903.8 506.74 L912.11 485.86 Z"
      /><path d="M912.11 485.86 L872.73 446.1 L840.16 473.4 L845.17 497.66 L903.8 506.74 L912.11 485.86 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M440 896.48 L432.29 904.38 L445.94 964.58 L456.77 966.23 L496.32 923.97 L496.15 923.11 L440 896.48 Z"
      /><path d="M440 896.48 L432.29 904.38 L445.94 964.58 L456.77 966.23 L496.32 923.97 L496.15 923.11 L440 896.48 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M1717.42 497.01 L1687.22 506.56 L1683.11 564.44 L1721.12 559.36 L1717.42 497.01 Z"
      /><path d="M1717.42 497.01 L1687.22 506.56 L1683.11 564.44 L1721.12 559.36 L1717.42 497.01 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M108.34 942.55 L105.46 946.86 L107.3 976.57 L154.41 996.65 L156.71 995.54 L172.22 969.16 L168.96 949.4 L108.34 942.55 Z"
      /><path d="M108.34 942.55 L105.46 946.86 L107.3 976.57 L154.41 996.65 L156.71 995.54 L172.22 969.16 L168.96 949.4 L108.34 942.55 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1610.45 998.31 L1629.38 1000.49 L1640.92 1016.11 L1634.17 1041.53 L1613.15 1052.92 L1586.51 1028.11 L1610.45 998.31 Z"
      /><path d="M1610.45 998.31 L1629.38 1000.49 L1640.92 1016.11 L1634.17 1041.53 L1613.15 1052.92 L1586.51 1028.11 L1610.45 998.31 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M749.06 275.39 L731.42 250.36 L699.26 253.72 L694.27 258.92 L700.68 290.37 L747.88 278.67 L749.06 275.39 Z"
      /><path d="M749.06 275.39 L731.42 250.36 L699.26 253.72 L694.27 258.92 L700.68 290.37 L747.88 278.67 L749.06 275.39 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1233.73 533.47 L1231.6801 561.6 L1205.77 570.4 L1181.79 545.07 L1197.17 517.92 L1213.23 513.76 L1233.73 533.47 Z"
      /><path d="M1233.73 533.47 L1231.6801 561.6 L1205.77 570.4 L1181.79 545.07 L1197.17 517.92 L1213.23 513.76 L1233.73 533.47 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M416.9 663.88 L398.99 621.76 L363.6 623.36 L352.01 635.46 L356.94 648.7 L393.6 673.26 L411.32 673.16 L416.9 663.88 Z"
      /><path d="M416.9 663.88 L398.99 621.76 L363.6 623.36 L352.01 635.46 L356.94 648.7 L393.6 673.26 L411.32 673.16 L416.9 663.88 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M135.54 1032.78 L99.7 1027.76 L84.25 1044.98 L88.1 1080 L141.2 1080 L145.1 1053.28 L135.54 1032.78 Z"
      /><path d="M135.54 1032.78 L99.7 1027.76 L84.25 1044.98 L88.1 1080 L141.2 1080 L145.1 1053.28 L135.54 1032.78 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1705.85 432.99 L1678.85 393.4 L1675.8 394.9 L1649.03 433.26 L1649.01 439 L1669.61 455.92 L1696.63 450.35 L1705.85 432.99 Z"
      /><path d="M1705.85 432.99 L1678.85 393.4 L1675.8 394.9 L1649.03 433.26 L1649.01 439 L1669.61 455.92 L1696.63 450.35 L1705.85 432.99 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1482.1 828.76 L1438.87 810.08 L1426 826.41 L1431.71 868.3 L1457.87 871.73 L1486.12 842.94 L1482.1 828.76 Z"
      /><path d="M1482.1 828.76 L1438.87 810.08 L1426 826.41 L1431.71 868.3 L1457.87 871.73 L1486.12 842.94 L1482.1 828.76 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1225.79 870.02 L1183.26 868.8 L1172.9301 878.74 L1178.9301 901.87 L1212.9399 913.57 L1226.24 907.47 L1227.04 871.53 L1225.79 870.02 Z"
      /><path d="M1225.79 870.02 L1183.26 868.8 L1172.9301 878.74 L1178.9301 901.87 L1212.9399 913.57 L1226.24 907.47 L1227.04 871.53 L1225.79 870.02 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M200.66 156.85 L228.02 160.6 L233.12 200.09 L191.62 216.34 L174.56 185.23 L200.66 156.85 Z"
      /><path d="M200.66 156.85 L228.02 160.6 L233.12 200.09 L191.62 216.34 L174.56 185.23 L200.66 156.85 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1261.96 994.31 L1262.95 996.09 L1260.28 1022.35 L1243.16 1038.62 L1230.4 1040.89 L1217.1801 1030.77 L1213.87 1013.05 L1237.03 985.87 L1261.96 994.31 Z"
      /><path d="M1261.96 994.31 L1262.95 996.09 L1260.28 1022.35 L1243.16 1038.62 L1230.4 1040.89 L1217.1801 1030.77 L1213.87 1013.05 L1237.03 985.87 L1261.96 994.31 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M515.88 941.16 L518.77 974.99 L483.66 994.61 L456.77 966.23 L496.32 923.97 L515.88 941.16 Z"
      /><path d="M515.88 941.16 L518.77 974.99 L483.66 994.61 L456.77 966.23 L496.32 923.97 L515.88 941.16 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1381.8199 277.55 L1325.02 265.41 L1315.33 271.52 L1324.33 307.61 L1359.61 316.26 L1383.7 280.18 L1381.8199 277.55 Z"
      /><path d="M1381.8199 277.55 L1325.02 265.41 L1315.33 271.52 L1324.33 307.61 L1359.61 316.26 L1383.7 280.18 L1381.8199 277.55 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1750.5 54.93 L1767.3199 72.9 L1753.01 118.95 L1752.36 119.35 L1713.0601 101.7 L1735.46 55.24 L1750.5 54.93 Z"
      /><path d="M1750.5 54.93 L1767.3199 72.9 L1753.01 118.95 L1752.36 119.35 L1713.0601 101.7 L1735.46 55.24 L1750.5 54.93 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M1477.99 642.06 L1489.5601 657.08 L1489.09 667.11 L1457.15 695.82 L1446.8199 693.29 L1428.92 662.82 L1433.1 642.15 L1477.99 642.06 Z"
      /><path d="M1477.99 642.06 L1489.5601 657.08 L1489.09 667.11 L1457.15 695.82 L1446.8199 693.29 L1428.92 662.82 L1433.1 642.15 L1477.99 642.06 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M482.72 447.92 L509.55 477.17 L490.43 502.02 L458.9 475.46 L462.49 460.86 L482.72 447.92 Z"
      /><path d="M482.72 447.92 L509.55 477.17 L490.43 502.02 L458.9 475.46 L462.49 460.86 L482.72 447.92 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1148.42 935.06 L1142.79 946.05 L1121.61 956.78 L1092.38 944.08 L1084.63 923.49 L1096.52 907.91 L1125.88 906.06 L1148.42 935.06 Z"
      /><path d="M1148.42 935.06 L1142.79 946.05 L1121.61 956.78 L1092.38 944.08 L1084.63 923.49 L1096.52 907.91 L1125.88 906.06 L1148.42 935.06 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M657.75 428.66 L645.17 426.9 L620.51 446.85 L628.91 476.75 L632.75 480.01 L671.49 474.05 L673.34 470.67 L657.75 428.66 Z"
      /><path d="M657.75 428.66 L645.17 426.9 L620.51 446.85 L628.91 476.75 L632.75 480.01 L671.49 474.05 L673.34 470.67 L657.75 428.66 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M445.52 55.89 L466.45 64 L469.53 70.69 L452.48 114.76 L418.48 107.99 L415.43 64.45 L445.52 55.89 Z"
      /><path d="M445.52 55.89 L466.45 64 L469.53 70.69 L452.48 114.76 L418.48 107.99 L415.43 64.45 L445.52 55.89 Z" style="fill:rgb(180,156,70); stroke:none;"
      /><path style="fill:none;" d="M769.07 1026.8101 L731.27 1031.6801 L728 1080 L775.5 1080 L769.07 1026.8101 Z"
      /><path d="M769.07 1026.8101 L731.27 1031.6801 L728 1080 L775.5 1080 L769.07 1026.8101 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M555.82 313.01 L524.92 308.38 L516.77 333.37 L542.7 359.3 L554.79 359.3 L555.82 313.01 Z"
      /><path d="M555.82 313.01 L524.92 308.38 L516.77 333.37 L542.7 359.3 L554.79 359.3 L555.82 313.01 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1183.85 830.15 L1183.26 868.8 L1172.9301 878.74 L1141.45 871.64 L1139.66 868.84 L1152.78 822.52 L1183.85 830.15 Z"
      /><path d="M1183.85 830.15 L1183.26 868.8 L1172.9301 878.74 L1141.45 871.64 L1139.66 868.84 L1152.78 822.52 L1183.85 830.15 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M669.14 610 L654.51 577.36 L626.12 578.99 L625.73 580.36 L636.09 612.09 L661.32 616.96 L669.14 610 Z"
      /><path d="M669.14 610 L654.51 577.36 L626.12 578.99 L625.73 580.36 L636.09 612.09 L661.32 616.96 L669.14 610 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1331.58 107.63 L1346.24 123.13 L1331.92 154.05 L1305.84 156.58 L1297.61 144.82 L1303.9301 110.89 L1331.58 107.63 Z"
      /><path d="M1331.58 107.63 L1346.24 123.13 L1331.92 154.05 L1305.84 156.58 L1297.61 144.82 L1303.9301 110.89 L1331.58 107.63 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1384.04 187.96 L1384.1899 224 L1378.5601 229.68 L1339.49 224.66 L1329.35 209.65 L1353.24 175.79 L1368.79 174.57 L1384.04 187.96 Z"
      /><path d="M1384.04 187.96 L1384.1899 224 L1378.5601 229.68 L1339.49 224.66 L1329.35 209.65 L1353.24 175.79 L1368.79 174.57 L1384.04 187.96 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M393.26 515.78 L433.22 528.29 L433.19 549.52 L402.82 573.21 L386.89 567.06 L379.05 526.24 L393.26 515.78 Z"
      /><path d="M393.26 515.78 L433.22 528.29 L433.19 549.52 L402.82 573.21 L386.89 567.06 L379.05 526.24 L393.26 515.78 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M307.49 703.68 L265.77 700.95 L253.38 725.63 L284.39 757.45 L286.21 757.11 L310.76 729.02 L307.49 703.68 Z"
      /><path d="M307.49 703.68 L265.77 700.95 L253.38 725.63 L284.39 757.45 L286.21 757.11 L310.76 729.02 L307.49 703.68 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M968.72 838.72 L932.61 839.71 L922.93 857.6 L925.76 866.67 L953.81 877.1 L974.68 852.69 L968.72 838.72 Z"
      /><path d="M968.72 838.72 L932.61 839.71 L922.93 857.6 L925.76 866.67 L953.81 877.1 L974.68 852.69 L968.72 838.72 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1860.7 183.37 L1840.87 166.19 L1802.0699 170.98 L1791.11 181.08 L1806.24 225.52 L1821.25 232.97 L1861.79 218.72 L1860.7 183.37 Z"
      /><path d="M1860.7 183.37 L1840.87 166.19 L1802.0699 170.98 L1791.11 181.08 L1806.24 225.52 L1821.25 232.97 L1861.79 218.72 L1860.7 183.37 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M736.25 598.88 L737.16 599.01 L759.06 637.67 L740.09 652.32 L704.99 646.62 L701.91 621.12 L736.25 598.88 Z"
      /><path d="M736.25 598.88 L737.16 599.01 L759.06 637.67 L740.09 652.32 L704.99 646.62 L701.91 621.12 L736.25 598.88 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M920.4 1029.73 L866.53 1022.19 L869.8 1080 L919.3 1080 L924.77 1034.8199 L920.4 1029.73 Z"
      /><path d="M920.4 1029.73 L866.53 1022.19 L869.8 1080 L919.3 1080 L924.77 1034.8199 L920.4 1029.73 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M96.83 534.46 L78.83 519.98 L61.35 546.95 L84 564.03 L90.45 560.05 L96.83 534.46 Z"
      /><path d="M96.83 534.46 L78.83 519.98 L61.35 546.95 L84 564.03 L90.45 560.05 L96.83 534.46 Z" style="fill:rgb(70,90,180); stroke:none;"
      /><path style="fill:none;" d="M530.38 131.69 L504.47 119.59 L480.4 131.57 L487.93 174.64 L516.66 170.99 L531.89 137.62 L530.38 131.69 Z"
      /><path d="M530.38 131.69 L504.47 119.59 L480.4 131.57 L487.93 174.64 L516.66 170.99 L531.89 137.62 L530.38 131.69 Z" style="fill:rgb(51,153,51); stroke:none;"
      /><path style="fill:none;" d="M1217.1801 1030.77 L1179 1048.79 L1181 1080 L1225 1080 L1230.4 1040.89 L1217.1801 1030.77 Z"
      /><path d="M1217.1801 1030.77 L1179 1048.79 L1181 1080 L1225 1080 L1230.4 1040.89 L1217.1801 1030.77 Z" style="fill:rgb(70,90,180); stroke:none;"
    /></g
  ></g
></svg
>
